-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity zm2_rom is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of zm2_rom is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"FF",x"FF",x"25",x"01",x"00",x"00",x"00",x"00", -- 0x0000
    x"50",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0010
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0020
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0030
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0040
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0050
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0060
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0070
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0080
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0088
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0090
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0100
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0110
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0120
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0130
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0140
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0150
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0170
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0180
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0190
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0210
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0260
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0280
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0290
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0300
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0310
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0320
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0330
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0340
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0350
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0360
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0370
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0380
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0390
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0400
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0410
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0420
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0430
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0440
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0450
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0458
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0460
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0468
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0470
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0480
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0490
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0540
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0548
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0550
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0560
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0570
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0580
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0588
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0590
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0610
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0618
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0620
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0630
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0638
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0640
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0648
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0650
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0658
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0660
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0668
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0670
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0678
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0680
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0688
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0690
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0698
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0700
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0710
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0720
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0730
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0740
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0750
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0760
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0770
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0780
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0798
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0800
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0810
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0818
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0820
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0828
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0830
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0838
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0840
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0848
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0850
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0858
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0860
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0868
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0870
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0878
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0880
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0890
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0898
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x08F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0900
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0908
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0910
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0918
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0920
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0928
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0930
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0938
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0940
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0948
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0950
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0958
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0960
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0968
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0970
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0978
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0980
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0988
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0990
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0998
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09A0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F08
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F20
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F28
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F48
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F50
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F78
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF8
    x"A0",x"04",x"B9",x"A0",x"F0",x"99",x"00",x"02", -- 0x1000
    x"88",x"10",x"F7",x"A2",x"FF",x"8E",x"20",x"02", -- 0x1008
    x"86",x"88",x"9A",x"A9",x"4C",x"85",x"A1",x"A2", -- 0x1010
    x"18",x"BD",x"A4",x"F0",x"95",x"BB",x"CA",x"D0", -- 0x1018
    x"F8",x"A2",x"12",x"BD",x"BD",x"F0",x"95",x"00", -- 0x1020
    x"CA",x"10",x"F8",x"A9",x"00",x"85",x"D8",x"85", -- 0x1028
    x"DB",x"85",x"B2",x"85",x"67",x"A9",x"0E",x"85", -- 0x1030
    x"64",x"A9",x"03",x"85",x"A0",x"A2",x"68",x"86", -- 0x1038
    x"65",x"A9",x"00",x"D0",x"1F",x"A0",x"00",x"E6", -- 0x1040
    x"11",x"D0",x"08",x"E6",x"12",x"A5",x"12",x"C9", -- 0x1048
    x"80",x"F0",x"1D",x"A9",x"55",x"91",x"11",x"D1", -- 0x1050
    x"11",x"D0",x"15",x"0A",x"91",x"11",x"D1",x"11", -- 0x1058
    x"F0",x"E5",x"D0",x"0C",x"20",x"50",x"E9",x"A5", -- 0x1060
    x"AC",x"C9",x"98",x"B0",x"B4",x"20",x"9E",x"E4", -- 0x1068
    x"A5",x"11",x"A4",x"12",x"C0",x"01",x"90",x"A9", -- 0x1070
    x"85",x"85",x"84",x"86",x"85",x"81",x"84",x"82", -- 0x1078
    x"A0",x"00",x"A2",x"04",x"84",x"79",x"86",x"7A", -- 0x1080
    x"98",x"91",x"79",x"E6",x"79",x"20",x"39",x"D8", -- 0x1088
    x"20",x"3F",x"D3",x"A5",x"85",x"38",x"E5",x"79", -- 0x1090
    x"AA",x"A5",x"86",x"E5",x"7A",x"20",x"2D",x"EA", -- 0x1098
    x"A9",x"DF",x"A0",x"F0",x"20",x"7A",x"D8",x"A9", -- 0x10A0
    x"49",x"A0",x"D1",x"85",x"01",x"84",x"02",x"6C", -- 0x10A8
    x"01",x"00",x"20",x"FC",x"D0",x"85",x"7F",x"84", -- 0x10B0
    x"80",x"38",x"A5",x"A6",x"E5",x"AA",x"A8",x"A5", -- 0x10B8
    x"A7",x"E5",x"AB",x"AA",x"E8",x"98",x"F0",x"24", -- 0x10C0
    x"38",x"49",x"FF",x"65",x"A6",x"85",x"A6",x"B0", -- 0x10C8
    x"03",x"C6",x"A7",x"38",x"98",x"49",x"FF",x"65", -- 0x10D0
    x"A4",x"85",x"A4",x"B0",x"08",x"C6",x"A5",x"90", -- 0x10D8
    x"04",x"B1",x"A6",x"91",x"A4",x"88",x"D0",x"F9", -- 0x10E0
    x"B1",x"A6",x"91",x"A4",x"C6",x"A7",x"C6",x"A5", -- 0x10E8
    x"CA",x"D0",x"F2",x"60",x"85",x"78",x"BA",x"E4", -- 0x10F0
    x"78",x"90",x"2E",x"60",x"C4",x"82",x"90",x"28", -- 0x10F8
    x"D0",x"04",x"C5",x"81",x"90",x"22",x"48",x"A2", -- 0x1100
    x"08",x"98",x"48",x"B5",x"A3",x"CA",x"10",x"FA", -- 0x1108
    x"20",x"86",x"E1",x"A2",x"F8",x"68",x"95",x"AC", -- 0x1110
    x"E8",x"30",x"FA",x"68",x"A8",x"68",x"C4",x"82", -- 0x1118
    x"90",x"06",x"D0",x"05",x"C5",x"81",x"B0",x"01", -- 0x1120
    x"60",x"A2",x"0C",x"20",x"39",x"D8",x"BD",x"47", -- 0x1128
    x"F6",x"BC",x"48",x"F6",x"20",x"7A",x"D8",x"20", -- 0x1130
    x"78",x"D3",x"A9",x"84",x"A0",x"F7",x"20",x"7A", -- 0x1138
    x"D8",x"A4",x"88",x"C8",x"F0",x"03",x"20",x"22", -- 0x1140
    x"EA",x"A9",x"00",x"85",x"DB",x"85",x"D8",x"A9", -- 0x1148
    x"95",x"A0",x"F7",x"20",x"7A",x"D8",x"20",x"3C", -- 0x1150
    x"D2",x"86",x"C3",x"84",x"C4",x"20",x"C2",x"00", -- 0x1158
    x"F0",x"F4",x"A2",x"FF",x"86",x"88",x"90",x"06", -- 0x1160
    x"20",x"6D",x"D2",x"4C",x"E2",x"D4",x"20",x"FA", -- 0x1168
    x"D6",x"20",x"6D",x"D2",x"84",x"5D",x"20",x"13", -- 0x1170
    x"D3",x"90",x"44",x"A0",x"01",x"B1",x"AA",x"85", -- 0x1178
    x"72",x"A5",x"7B",x"85",x"71",x"A5",x"AB",x"85", -- 0x1180
    x"74",x"A5",x"AA",x"88",x"F1",x"AA",x"18",x"65", -- 0x1188
    x"7B",x"85",x"7B",x"85",x"73",x"A5",x"7C",x"69", -- 0x1190
    x"FF",x"85",x"7C",x"E5",x"AB",x"AA",x"38",x"A5", -- 0x1198
    x"AA",x"E5",x"7B",x"A8",x"B0",x"03",x"E8",x"C6", -- 0x11A0
    x"74",x"18",x"65",x"71",x"90",x"03",x"C6",x"72", -- 0x11A8
    x"18",x"B1",x"71",x"91",x"73",x"C8",x"D0",x"F9", -- 0x11B0
    x"E6",x"72",x"E6",x"74",x"CA",x"D0",x"F2",x"AD", -- 0x11B8
    x"21",x"02",x"F0",x"3F",x"A5",x"85",x"A4",x"86", -- 0x11C0
    x"85",x"81",x"84",x"82",x"A5",x"7B",x"85",x"A6", -- 0x11C8
    x"A4",x"7C",x"84",x"A7",x"65",x"5D",x"90",x"01", -- 0x11D0
    x"C8",x"85",x"A4",x"84",x"A5",x"20",x"B2",x"D0", -- 0x11D8
    x"A5",x"7F",x"A4",x"80",x"85",x"7B",x"84",x"7C", -- 0x11E0
    x"A4",x"5D",x"88",x"B9",x"1D",x"02",x"91",x"AA", -- 0x11E8
    x"88",x"C0",x"03",x"D0",x"F6",x"A5",x"12",x"91", -- 0x11F0
    x"AA",x"88",x"A5",x"11",x"91",x"AA",x"88",x"A9", -- 0x11F8
    x"FF",x"91",x"AA",x"20",x"54",x"D3",x"A6",x"79", -- 0x1200
    x"A5",x"7A",x"A0",x"01",x"86",x"71",x"85",x"72", -- 0x1208
    x"B1",x"71",x"F0",x"18",x"A0",x"04",x"C8",x"B1", -- 0x1210
    x"71",x"D0",x"FB",x"38",x"98",x"65",x"71",x"AA", -- 0x1218
    x"A0",x"00",x"91",x"71",x"98",x"65",x"72",x"C8", -- 0x1220
    x"91",x"71",x"90",x"E0",x"4C",x"56",x"D1",x"20", -- 0x1228
    x"92",x"D8",x"20",x"8F",x"D8",x"D0",x"05",x"20", -- 0x1230
    x"94",x"D8",x"CA",x"2C",x"A2",x"00",x"20",x"94", -- 0x1238
    x"F0",x"90",x"FB",x"F0",x"F9",x"C9",x"07",x"F0", -- 0x1240
    x"10",x"C9",x"0D",x"F0",x"19",x"E0",x"00",x"D0", -- 0x1248
    x"04",x"C9",x"21",x"90",x"E9",x"C9",x"08",x"F0", -- 0x1250
    x"DE",x"E0",x"47",x"B0",x"0C",x"9D",x"21",x"02", -- 0x1258
    x"E8",x"20",x"94",x"D8",x"D0",x"D8",x"4C",x"30", -- 0x1260
    x"D8",x"A9",x"07",x"D0",x"F4",x"A0",x"FF",x"38", -- 0x1268
    x"A5",x"C3",x"E9",x"21",x"AA",x"86",x"60",x"BD", -- 0x1270
    x"21",x"02",x"F0",x"51",x"C9",x"5F",x"B0",x"4D", -- 0x1278
    x"C9",x"3C",x"B0",x"0E",x"C9",x"30",x"B0",x"45", -- 0x1280
    x"85",x"5C",x"C9",x"22",x"F0",x"61",x"C9",x"2A", -- 0x1288
    x"90",x"3B",x"24",x"60",x"70",x"37",x"86",x"78", -- 0x1290
    x"84",x"BA",x"A0",x"B6",x"84",x"73",x"A0",x"F2", -- 0x1298
    x"84",x"74",x"A0",x"00",x"D1",x"73",x"F0",x"05", -- 0x12A0
    x"90",x"21",x"C8",x"D0",x"F7",x"98",x"0A",x"AA", -- 0x12A8
    x"BD",x"D4",x"F2",x"85",x"73",x"BD",x"D5",x"F2", -- 0x12B0
    x"85",x"74",x"A0",x"FF",x"A6",x"78",x"C8",x"B1", -- 0x12B8
    x"73",x"30",x"08",x"E8",x"DD",x"21",x"02",x"F0", -- 0x12C0
    x"F5",x"D0",x"2B",x"A4",x"BA",x"E8",x"C8",x"99", -- 0x12C8
    x"21",x"02",x"C9",x"00",x"F0",x"32",x"E9",x"3A", -- 0x12D0
    x"F0",x"04",x"C9",x"49",x"D0",x"02",x"85",x"60", -- 0x12D8
    x"49",x"57",x"D0",x"93",x"85",x"5C",x"BD",x"21", -- 0x12E0
    x"02",x"F0",x"E2",x"C5",x"5C",x"F0",x"DE",x"C8", -- 0x12E8
    x"99",x"21",x"02",x"E8",x"D0",x"F0",x"A6",x"78", -- 0x12F0
    x"B1",x"73",x"08",x"C8",x"28",x"10",x"F9",x"B1", -- 0x12F8
    x"73",x"D0",x"BE",x"BD",x"21",x"02",x"10",x"C3", -- 0x1300
    x"C8",x"C8",x"99",x"21",x"02",x"C8",x"C8",x"C8", -- 0x1308
    x"C6",x"C3",x"60",x"A5",x"79",x"A6",x"7A",x"A0", -- 0x1310
    x"01",x"85",x"AA",x"86",x"AB",x"B1",x"AA",x"F0", -- 0x1318
    x"1A",x"A0",x"03",x"B1",x"AA",x"88",x"C5",x"12", -- 0x1320
    x"D0",x"04",x"B1",x"AA",x"C5",x"11",x"B0",x"09", -- 0x1328
    x"88",x"B1",x"AA",x"AA",x"88",x"B1",x"AA",x"90", -- 0x1330
    x"DE",x"F0",x"01",x"18",x"60",x"D0",x"FD",x"A9", -- 0x1338
    x"00",x"A8",x"91",x"79",x"C8",x"91",x"79",x"18", -- 0x1340
    x"A5",x"79",x"69",x"02",x"85",x"7B",x"A5",x"7A", -- 0x1348
    x"69",x"00",x"85",x"7C",x"18",x"A5",x"79",x"69", -- 0x1350
    x"FF",x"85",x"C3",x"A5",x"7A",x"69",x"FF",x"85", -- 0x1358
    x"C4",x"A5",x"85",x"A4",x"86",x"85",x"81",x"84", -- 0x1360
    x"82",x"A5",x"7B",x"A4",x"7C",x"85",x"7D",x"84", -- 0x1368
    x"7E",x"85",x"7F",x"84",x"80",x"20",x"33",x"D5", -- 0x1370
    x"A2",x"68",x"86",x"65",x"68",x"AA",x"68",x"8E", -- 0x1378
    x"FE",x"01",x"8D",x"FF",x"01",x"A2",x"FD",x"9A", -- 0x1380
    x"A9",x"00",x"85",x"8C",x"85",x"61",x"60",x"F0", -- 0x1388
    x"D0",x"60",x"90",x"06",x"F0",x"04",x"C9",x"B6", -- 0x1390
    x"D0",x"F4",x"20",x"FA",x"D6",x"20",x"13",x"D3", -- 0x1398
    x"20",x"C2",x"00",x"F0",x"0C",x"C9",x"B6",x"D0", -- 0x13A0
    x"93",x"20",x"BC",x"00",x"20",x"FA",x"D6",x"D0", -- 0x13A8
    x"8B",x"A5",x"11",x"05",x"12",x"D0",x"06",x"A9", -- 0x13B0
    x"FF",x"85",x"11",x"85",x"12",x"A0",x"01",x"84", -- 0x13B8
    x"60",x"20",x"39",x"D8",x"B1",x"AA",x"F0",x"3E", -- 0x13C0
    x"20",x"03",x"D5",x"C8",x"B1",x"AA",x"AA",x"C8", -- 0x13C8
    x"B1",x"AA",x"C5",x"12",x"D0",x"04",x"E4",x"11", -- 0x13D0
    x"F0",x"02",x"B0",x"2A",x"84",x"97",x"20",x"2D", -- 0x13D8
    x"EA",x"A9",x"20",x"A4",x"97",x"29",x"7F",x"20", -- 0x13E0
    x"94",x"D8",x"C9",x"22",x"D0",x"06",x"A5",x"60", -- 0x13E8
    x"49",x"FF",x"85",x"60",x"C8",x"B1",x"AA",x"D0", -- 0x13F0
    x"0E",x"A8",x"B1",x"AA",x"AA",x"C8",x"B1",x"AA", -- 0x13F8
    x"86",x"AA",x"85",x"AB",x"D0",x"B7",x"60",x"10", -- 0x1400
    x"DE",x"24",x"60",x"30",x"DA",x"A2",x"F4",x"0A", -- 0x1408
    x"0A",x"90",x"02",x"E8",x"18",x"69",x"B3",x"90", -- 0x1410
    x"01",x"E8",x"85",x"73",x"86",x"74",x"84",x"97", -- 0x1418
    x"A0",x"00",x"B1",x"73",x"AA",x"C8",x"B1",x"73", -- 0x1420
    x"CA",x"F0",x"B8",x"20",x"94",x"D8",x"C8",x"B1", -- 0x1428
    x"73",x"48",x"C8",x"B1",x"73",x"A0",x"00",x"85", -- 0x1430
    x"74",x"68",x"85",x"73",x"B1",x"73",x"CA",x"F0", -- 0x1438
    x"A2",x"20",x"94",x"D8",x"C8",x"D0",x"F5",x"A9", -- 0x1440
    x"80",x"85",x"61",x"20",x"59",x"D7",x"68",x"68", -- 0x1448
    x"A9",x"10",x"20",x"F4",x"D0",x"20",x"8C",x"D6", -- 0x1450
    x"18",x"98",x"65",x"C3",x"48",x"A5",x"C4",x"69", -- 0x1458
    x"00",x"48",x"A5",x"88",x"48",x"A5",x"87",x"48", -- 0x1460
    x"A9",x"AC",x"20",x"98",x"DB",x"20",x"77",x"DA", -- 0x1468
    x"20",x"74",x"DA",x"A5",x"B0",x"09",x"7F",x"25", -- 0x1470
    x"AD",x"85",x"AD",x"A9",x"86",x"A0",x"D4",x"85", -- 0x1478
    x"71",x"84",x"72",x"4C",x"2B",x"DB",x"A9",x"86", -- 0x1480
    x"A0",x"F1",x"20",x"27",x"E8",x"20",x"C2",x"00", -- 0x1488
    x"C9",x"B1",x"D0",x"06",x"20",x"BC",x"00",x"20", -- 0x1490
    x"74",x"DA",x"20",x"93",x"E8",x"85",x"B0",x"20", -- 0x1498
    x"20",x"DB",x"A5",x"98",x"48",x"A5",x"97",x"48", -- 0x14A0
    x"A9",x"81",x"48",x"20",x"03",x"D5",x"A5",x"C3", -- 0x14A8
    x"A4",x"C4",x"A6",x"88",x"E8",x"F0",x"04",x"85", -- 0x14B0
    x"8B",x"84",x"8C",x"A0",x"00",x"B1",x"C3",x"F0", -- 0x14B8
    x"07",x"C9",x"3A",x"F0",x"1D",x"4C",x"A9",x"DB", -- 0x14C0
    x"A0",x"02",x"B1",x"C3",x"18",x"F0",x"56",x"C8", -- 0x14C8
    x"B1",x"C3",x"85",x"87",x"C8",x"B1",x"C3",x"85", -- 0x14D0
    x"88",x"98",x"65",x"C3",x"85",x"C3",x"90",x"02", -- 0x14D8
    x"E6",x"C4",x"20",x"BC",x"00",x"20",x"EB",x"D4", -- 0x14E0
    x"4C",x"AB",x"D4",x"F0",x"54",x"0A",x"B0",x"03", -- 0x14E8
    x"4C",x"59",x"D7",x"C9",x"56",x"B0",x"CE",x"A8", -- 0x14F0
    x"B9",x"AE",x"F1",x"48",x"B9",x"AD",x"F1",x"48", -- 0x14F8
    x"4C",x"BC",x"00",x"6C",x"03",x"02",x"C9",x"03", -- 0x1500
    x"B0",x"01",x"18",x"D0",x"67",x"A5",x"C4",x"49", -- 0x1508
    x"02",x"F0",x"10",x"49",x"02",x"A4",x"C3",x"84", -- 0x1510
    x"8B",x"85",x"8C",x"A5",x"87",x"A4",x"88",x"85", -- 0x1518
    x"89",x"84",x"8A",x"68",x"68",x"90",x"07",x"A9", -- 0x1520
    x"7C",x"A0",x"F7",x"4C",x"3E",x"D1",x"4C",x"49", -- 0x1528
    x"D1",x"D0",x"0F",x"38",x"A5",x"79",x"E9",x"01", -- 0x1530
    x"A4",x"7A",x"B0",x"01",x"88",x"85",x"8F",x"84", -- 0x1538
    x"90",x"60",x"20",x"FA",x"D6",x"20",x"8F",x"D6", -- 0x1540
    x"A5",x"88",x"C5",x"12",x"B0",x"0B",x"98",x"38", -- 0x1548
    x"65",x"C3",x"A6",x"C4",x"90",x"07",x"E8",x"B0", -- 0x1550
    x"04",x"A5",x"79",x"A6",x"7A",x"20",x"17",x"D3", -- 0x1558
    x"B0",x"03",x"4C",x"61",x"D6",x"A5",x"AA",x"E9", -- 0x1560
    x"01",x"A4",x"AB",x"B0",x"D0",x"90",x"CD",x"20", -- 0x1568
    x"33",x"E4",x"86",x"0D",x"60",x"D0",x"FD",x"A4", -- 0x1570
    x"8C",x"D0",x"05",x"A2",x"1E",x"4C",x"2B",x"D1", -- 0x1578
    x"A9",x"93",x"20",x"BE",x"EE",x"A9",x"93",x"20", -- 0x1580
    x"C1",x"EE",x"84",x"C4",x"A5",x"8B",x"85",x"C3", -- 0x1588
    x"A5",x"89",x"A4",x"8A",x"85",x"87",x"84",x"88", -- 0x1590
    x"60",x"D0",x"03",x"4C",x"54",x"D3",x"20",x"61", -- 0x1598
    x"D3",x"F0",x"2E",x"A9",x"05",x"20",x"F4",x"D0", -- 0x15A0
    x"A5",x"C4",x"48",x"A5",x"C3",x"48",x"A5",x"88", -- 0x15A8
    x"48",x"A5",x"87",x"48",x"A9",x"9D",x"48",x"20", -- 0x15B0
    x"C2",x"00",x"4C",x"AB",x"D4",x"A9",x"05",x"20", -- 0x15B8
    x"F4",x"D0",x"A5",x"C4",x"48",x"A5",x"C3",x"48", -- 0x15C0
    x"A5",x"88",x"48",x"A5",x"87",x"48",x"A9",x"8D", -- 0x15C8
    x"48",x"20",x"C2",x"00",x"20",x"DA",x"D5",x"4C", -- 0x15D0
    x"AB",x"D4",x"20",x"FA",x"D6",x"20",x"8F",x"D6", -- 0x15D8
    x"A5",x"88",x"C5",x"12",x"B0",x"0B",x"98",x"38", -- 0x15E0
    x"65",x"C3",x"A6",x"C4",x"90",x"07",x"E8",x"B0", -- 0x15E8
    x"04",x"A5",x"79",x"A6",x"7A",x"20",x"17",x"D3", -- 0x15F0
    x"90",x"67",x"A5",x"AA",x"E9",x"01",x"85",x"C3", -- 0x15F8
    x"A5",x"AB",x"E9",x"00",x"85",x"C4",x"60",x"A2", -- 0x1600
    x"22",x"4C",x"2B",x"D1",x"A8",x"BA",x"BD",x"03", -- 0x1608
    x"01",x"C9",x"9D",x"D0",x"F2",x"E8",x"E8",x"9A", -- 0x1610
    x"98",x"F0",x"20",x"C9",x"3A",x"F0",x"1C",x"E9", -- 0x1618
    x"B2",x"AA",x"F0",x"04",x"CA",x"D0",x"62",x"CA", -- 0x1620
    x"86",x"98",x"20",x"BC",x"00",x"20",x"88",x"DA", -- 0x1628
    x"A5",x"AC",x"F0",x"02",x"A9",x"FF",x"BA",x"45", -- 0x1630
    x"98",x"D0",x"1A",x"BD",x"02",x"01",x"85",x"87", -- 0x1638
    x"BD",x"03",x"01",x"85",x"88",x"BD",x"04",x"01", -- 0x1640
    x"85",x"C3",x"BD",x"05",x"01",x"85",x"C4",x"20", -- 0x1648
    x"C2",x"00",x"4C",x"AB",x"D4",x"E8",x"E8",x"E8", -- 0x1650
    x"E8",x"E8",x"9A",x"4C",x"7B",x"D6",x"A2",x"04", -- 0x1658
    x"2C",x"A2",x"0E",x"4C",x"2B",x"D1",x"D0",x"9E", -- 0x1660
    x"68",x"68",x"68",x"C9",x"8D",x"D0",x"EF",x"68", -- 0x1668
    x"85",x"87",x"68",x"85",x"88",x"68",x"85",x"C3", -- 0x1670
    x"68",x"85",x"C4",x"20",x"8C",x"D6",x"98",x"18", -- 0x1678
    x"65",x"C3",x"85",x"C3",x"90",x"02",x"E6",x"C4", -- 0x1680
    x"60",x"4C",x"A9",x"DB",x"A2",x"3A",x"2C",x"A2", -- 0x1688
    x"00",x"A0",x"00",x"84",x"5C",x"8A",x"45",x"5C", -- 0x1690
    x"85",x"5C",x"B1",x"C3",x"F0",x"EA",x"C5",x"5C", -- 0x1698
    x"F0",x"E6",x"C8",x"C9",x"22",x"D0",x"F3",x"F0", -- 0x16A0
    x"EC",x"20",x"88",x"DA",x"20",x"C2",x"00",x"C9", -- 0x16A8
    x"89",x"F0",x"05",x"A9",x"AF",x"20",x"98",x"DB", -- 0x16B0
    x"A5",x"AC",x"D0",x"05",x"20",x"8F",x"D6",x"F0", -- 0x16B8
    x"BD",x"20",x"C2",x"00",x"B0",x"03",x"4C",x"DA", -- 0x16C0
    x"D5",x"4C",x"EB",x"D4",x"C9",x"A9",x"D0",x"03", -- 0x16C8
    x"4C",x"E2",x"EE",x"C9",x"AA",x"D0",x"03",x"4C", -- 0x16D0
    x"E6",x"EE",x"20",x"33",x"E4",x"48",x"C9",x"8D", -- 0x16D8
    x"F0",x"04",x"C9",x"89",x"D0",x"A3",x"C6",x"AF", -- 0x16E0
    x"D0",x"04",x"68",x"4C",x"ED",x"D4",x"20",x"BC", -- 0x16E8
    x"00",x"20",x"FA",x"D6",x"C9",x"2C",x"F0",x"EE", -- 0x16F0
    x"68",x"60",x"A2",x"00",x"86",x"11",x"86",x"12", -- 0x16F8
    x"B0",x"F7",x"E0",x"19",x"A8",x"B0",x"DD",x"E9", -- 0x1700
    x"2F",x"A8",x"A5",x"11",x"0A",x"26",x"12",x"0A", -- 0x1708
    x"26",x"12",x"65",x"11",x"85",x"11",x"8A",x"65", -- 0x1710
    x"12",x"06",x"11",x"2A",x"AA",x"98",x"65",x"11", -- 0x1718
    x"85",x"11",x"90",x"01",x"E8",x"20",x"BC",x"00", -- 0x1720
    x"4C",x"FE",x"D6",x"A9",x"8A",x"2C",x"A9",x"86", -- 0x1728
    x"48",x"20",x"51",x"DD",x"A6",x"5F",x"30",x"1E", -- 0x1730
    x"85",x"97",x"84",x"98",x"20",x"27",x"E8",x"68", -- 0x1738
    x"48",x"A0",x"F1",x"20",x"65",x"E5",x"20",x"4D", -- 0x1740
    x"E8",x"20",x"C2",x"00",x"C9",x"2C",x"D0",x"A8", -- 0x1748
    x"20",x"BC",x"00",x"4C",x"31",x"D7",x"4C",x"83", -- 0x1750
    x"DA",x"20",x"51",x"DD",x"85",x"97",x"84",x"98", -- 0x1758
    x"A9",x"C0",x"20",x"98",x"DB",x"A5",x"5F",x"48", -- 0x1760
    x"20",x"88",x"DA",x"68",x"2A",x"20",x"7A",x"DA", -- 0x1768
    x"D0",x"03",x"4C",x"4D",x"E8",x"A0",x"02",x"B1", -- 0x1770
    x"AE",x"C5",x"82",x"90",x"17",x"D0",x"07",x"88", -- 0x1778
    x"B1",x"AE",x"C5",x"81",x"90",x"0E",x"A4",x"AF", -- 0x1780
    x"C4",x"7C",x"90",x"08",x"D0",x"0D",x"A5",x"AE", -- 0x1788
    x"C5",x"7B",x"B0",x"07",x"A5",x"AE",x"A4",x"AF", -- 0x1790
    x"4C",x"B1",x"D7",x"A0",x"00",x"B1",x"AE",x"20", -- 0x1798
    x"D9",x"E0",x"A5",x"9E",x"A4",x"9F",x"85",x"B8", -- 0x17A0
    x"84",x"B9",x"20",x"B8",x"E2",x"A9",x"AC",x"A0", -- 0x17A8
    x"00",x"85",x"9E",x"84",x"9F",x"20",x"1A",x"E3", -- 0x17B0
    x"A0",x"00",x"B1",x"9E",x"91",x"97",x"C8",x"B1", -- 0x17B8
    x"9E",x"91",x"97",x"C8",x"B1",x"9E",x"91",x"97", -- 0x17C0
    x"60",x"20",x"51",x"DD",x"85",x"97",x"84",x"98", -- 0x17C8
    x"20",x"AA",x"EE",x"A6",x"5F",x"30",x"07",x"A8", -- 0x17D0
    x"20",x"0D",x"E0",x"4C",x"4D",x"E8",x"48",x"A9", -- 0x17D8
    x"01",x"B0",x"01",x"68",x"20",x"E1",x"E0",x"F0", -- 0x17E0
    x"05",x"68",x"A0",x"00",x"91",x"AD",x"20",x"2C", -- 0x17E8
    x"E1",x"4C",x"75",x"D7",x"20",x"7D",x"D8",x"20", -- 0x17F0
    x"C2",x"00",x"F0",x"3D",x"F0",x"CA",x"C9",x"AB", -- 0x17F8
    x"F0",x"56",x"C9",x"AE",x"F0",x"52",x"C9",x"2C", -- 0x1800
    x"F0",x"38",x"C9",x"3B",x"F0",x"66",x"20",x"88", -- 0x1808
    x"DA",x"24",x"5F",x"30",x"DF",x"20",x"40",x"EA", -- 0x1810
    x"20",x"EB",x"E0",x"A0",x"00",x"A5",x"0F",x"F0", -- 0x1818
    x"0A",x"38",x"E5",x"0E",x"F1",x"AE",x"B0",x"03", -- 0x1820
    x"20",x"39",x"D8",x"20",x"7D",x"D8",x"F0",x"C7", -- 0x1828
    x"A9",x"00",x"9D",x"21",x"02",x"A2",x"21",x"A0", -- 0x1830
    x"02",x"A9",x"0D",x"20",x"94",x"D8",x"A9",x"0A", -- 0x1838
    x"D0",x"52",x"A5",x"0E",x"C5",x"10",x"90",x"05", -- 0x1840
    x"20",x"39",x"D8",x"D0",x"27",x"38",x"E5",x"64", -- 0x1848
    x"B0",x"FC",x"49",x"FF",x"69",x"01",x"D0",x"12", -- 0x1850
    x"48",x"20",x"30",x"E4",x"C9",x"29",x"D0",x"7B", -- 0x1858
    x"68",x"C9",x"AB",x"D0",x"06",x"8A",x"E5",x"0E", -- 0x1860
    x"90",x"0A",x"AA",x"8A",x"F0",x"06",x"20",x"8F", -- 0x1868
    x"D8",x"CA",x"D0",x"FA",x"20",x"BC",x"00",x"4C", -- 0x1870
    x"FC",x"D7",x"20",x"EB",x"E0",x"20",x"E5",x"E2", -- 0x1878
    x"A0",x"00",x"AA",x"F0",x"49",x"B1",x"71",x"20", -- 0x1880
    x"94",x"D8",x"C8",x"CA",x"D0",x"F7",x"60",x"A9", -- 0x1888
    x"20",x"2C",x"A9",x"3F",x"C9",x"20",x"90",x"19", -- 0x1890
    x"48",x"A5",x"0F",x"D0",x"0A",x"A5",x"0E",x"E5", -- 0x1898
    x"64",x"D0",x"0B",x"85",x"0E",x"F0",x"07",x"C5", -- 0x18A0
    x"0E",x"D0",x"03",x"20",x"39",x"D8",x"E6",x"0E", -- 0x18A8
    x"68",x"20",x"97",x"F0",x"C9",x"0D",x"D0",x"14", -- 0x18B0
    x"86",x"78",x"A6",x"0D",x"F0",x"0A",x"A9",x"00", -- 0x18B8
    x"20",x"94",x"D8",x"CA",x"D0",x"FA",x"A9",x"0D", -- 0x18C0
    x"86",x"0E",x"A6",x"78",x"29",x"FF",x"60",x"A5", -- 0x18C8
    x"62",x"10",x"0B",x"A5",x"8D",x"A4",x"8E",x"85", -- 0x18D0
    x"87",x"84",x"88",x"4C",x"A9",x"DB",x"A9",x"B0", -- 0x18D8
    x"A0",x"F7",x"20",x"7A",x"D8",x"A5",x"8B",x"A4", -- 0x18E0
    x"8C",x"85",x"C3",x"84",x"C4",x"60",x"C9",x"22", -- 0x18E8
    x"D0",x"0B",x"20",x"65",x"DB",x"A9",x"3B",x"20", -- 0x18F0
    x"98",x"DB",x"20",x"7D",x"D8",x"20",x"11",x"E0", -- 0x18F8
    x"20",x"2F",x"D2",x"A9",x"00",x"CD",x"21",x"02", -- 0x1900
    x"D0",x"0A",x"18",x"4C",x"1B",x"D5",x"A6",x"8F", -- 0x1908
    x"A4",x"90",x"A9",x"80",x"85",x"62",x"86",x"91", -- 0x1910
    x"84",x"92",x"20",x"51",x"DD",x"85",x"97",x"84", -- 0x1918
    x"98",x"A5",x"C3",x"A4",x"C4",x"85",x"11",x"84", -- 0x1920
    x"12",x"A6",x"91",x"A4",x"92",x"86",x"C3",x"84", -- 0x1928
    x"C4",x"20",x"C2",x"00",x"D0",x"11",x"24",x"62", -- 0x1930
    x"30",x"65",x"20",x"92",x"D8",x"20",x"2F",x"D2", -- 0x1938
    x"86",x"C3",x"84",x"C4",x"20",x"C2",x"00",x"24", -- 0x1940
    x"5F",x"10",x"24",x"85",x"5B",x"C9",x"22",x"F0", -- 0x1948
    x"07",x"A9",x"3A",x"85",x"5B",x"A9",x"2C",x"18", -- 0x1950
    x"85",x"5C",x"A5",x"C3",x"A4",x"C4",x"69",x"00", -- 0x1958
    x"90",x"01",x"C8",x"20",x"F1",x"E0",x"20",x"76", -- 0x1960
    x"E4",x"20",x"75",x"D7",x"4C",x"75",x"D9",x"20", -- 0x1968
    x"50",x"E9",x"20",x"4D",x"E8",x"20",x"C2",x"00", -- 0x1970
    x"F0",x"0A",x"C9",x"2C",x"F0",x"03",x"4C",x"CF", -- 0x1978
    x"D8",x"20",x"BC",x"00",x"A5",x"C3",x"A4",x"C4", -- 0x1980
    x"85",x"91",x"84",x"92",x"A5",x"11",x"A4",x"12", -- 0x1988
    x"85",x"C3",x"84",x"C4",x"20",x"C2",x"00",x"F0", -- 0x1990
    x"2C",x"20",x"A5",x"DB",x"4C",x"1A",x"D9",x"20", -- 0x1998
    x"8C",x"D6",x"C8",x"AA",x"D0",x"12",x"A2",x"06", -- 0x19A0
    x"C8",x"B1",x"C3",x"F0",x"73",x"C8",x"B1",x"C3", -- 0x19A8
    x"85",x"8D",x"C8",x"B1",x"C3",x"C8",x"85",x"8E", -- 0x19B0
    x"B1",x"C3",x"C8",x"AA",x"20",x"7E",x"D6",x"E0", -- 0x19B8
    x"83",x"F0",x"81",x"D0",x"DA",x"A5",x"91",x"A4", -- 0x19C0
    x"92",x"A6",x"62",x"10",x"03",x"4C",x"3D",x"D5", -- 0x19C8
    x"A0",x"00",x"B1",x"91",x"D0",x"01",x"60",x"A9", -- 0x19D0
    x"9F",x"A0",x"F7",x"4C",x"7A",x"D8",x"BA",x"E8", -- 0x19D8
    x"E8",x"E8",x"E8",x"BD",x"01",x"01",x"C9",x"81", -- 0x19E0
    x"D0",x"21",x"A5",x"98",x"D0",x"0A",x"BD",x"02", -- 0x19E8
    x"01",x"85",x"97",x"BD",x"03",x"01",x"85",x"98", -- 0x19F0
    x"DD",x"03",x"01",x"D0",x"07",x"A5",x"97",x"DD", -- 0x19F8
    x"02",x"01",x"F0",x"07",x"8A",x"18",x"69",x"10", -- 0x1A00
    x"AA",x"D0",x"D8",x"60",x"D0",x"04",x"A0",x"00", -- 0x1A08
    x"F0",x"03",x"20",x"51",x"DD",x"85",x"97",x"84", -- 0x1A10
    x"98",x"20",x"DE",x"D9",x"F0",x"04",x"A2",x"00", -- 0x1A18
    x"F0",x"63",x"9A",x"8A",x"38",x"E9",x"F7",x"85", -- 0x1A20
    x"73",x"69",x"FB",x"A0",x"01",x"20",x"27",x"E8", -- 0x1A28
    x"BA",x"BD",x"08",x"01",x"85",x"B0",x"A5",x"97", -- 0x1A30
    x"A4",x"98",x"20",x"65",x"E5",x"20",x"4D",x"E8", -- 0x1A38
    x"A0",x"01",x"20",x"C3",x"E8",x"BA",x"DD",x"08", -- 0x1A40
    x"01",x"F0",x"17",x"BD",x"0D",x"01",x"85",x"87", -- 0x1A48
    x"BD",x"0E",x"01",x"85",x"88",x"BD",x"10",x"01", -- 0x1A50
    x"85",x"C3",x"BD",x"0F",x"01",x"85",x"C4",x"4C", -- 0x1A58
    x"AB",x"D4",x"8A",x"69",x"0F",x"AA",x"9A",x"20", -- 0x1A60
    x"C2",x"00",x"C9",x"2C",x"D0",x"F1",x"20",x"BC", -- 0x1A68
    x"00",x"20",x"12",x"DA",x"20",x"88",x"DA",x"18", -- 0x1A70
    x"24",x"38",x"24",x"5F",x"30",x"03",x"B0",x"03", -- 0x1A78
    x"60",x"B0",x"FD",x"A2",x"18",x"4C",x"2B",x"D1", -- 0x1A80
    x"A6",x"C3",x"D0",x"02",x"C6",x"C4",x"C6",x"C3", -- 0x1A88
    x"A9",x"00",x"48",x"A9",x"02",x"20",x"F4",x"D0", -- 0x1A90
    x"20",x"74",x"DB",x"A9",x"00",x"85",x"9B",x"20", -- 0x1A98
    x"C2",x"00",x"38",x"E9",x"BF",x"90",x"17",x"C9", -- 0x1AA0
    x"03",x"B0",x"13",x"C9",x"01",x"2A",x"49",x"01", -- 0x1AA8
    x"45",x"9B",x"C5",x"9B",x"90",x"67",x"85",x"9B", -- 0x1AB0
    x"20",x"BC",x"00",x"4C",x"A2",x"DA",x"A6",x"9B", -- 0x1AB8
    x"D0",x"2C",x"B0",x"79",x"69",x"0A",x"90",x"75", -- 0x1AC0
    x"D0",x"07",x"24",x"5F",x"10",x"03",x"4C",x"7B", -- 0x1AC8
    x"E2",x"85",x"71",x"0A",x"65",x"71",x"A8",x"68", -- 0x1AD0
    x"D9",x"8F",x"F2",x"B0",x"65",x"20",x"77",x"DA", -- 0x1AD8
    x"48",x"20",x"09",x"DB",x"68",x"A4",x"99",x"10", -- 0x1AE0
    x"19",x"AA",x"F0",x"76",x"D0",x"5D",x"26",x"5F", -- 0x1AE8
    x"8A",x"85",x"5F",x"2A",x"A6",x"C3",x"D0",x"02", -- 0x1AF0
    x"C6",x"C4",x"C6",x"C3",x"A0",x"24",x"85",x"9B", -- 0x1AF8
    x"D0",x"D5",x"D9",x"8F",x"F2",x"B0",x"44",x"90", -- 0x1B00
    x"D7",x"B9",x"91",x"F2",x"48",x"B9",x"90",x"F2", -- 0x1B08
    x"48",x"20",x"20",x"DB",x"A5",x"9B",x"48",x"B9", -- 0x1B10
    x"8F",x"F2",x"4C",x"92",x"DA",x"4C",x"A9",x"DB", -- 0x1B18
    x"68",x"85",x"71",x"E6",x"71",x"68",x"85",x"72", -- 0x1B20
    x"A5",x"B0",x"48",x"20",x"83",x"E8",x"A5",x"AF", -- 0x1B28
    x"48",x"A5",x"AE",x"48",x"A5",x"AD",x"48",x"A5", -- 0x1B30
    x"AC",x"48",x"6C",x"71",x"00",x"A0",x"FF",x"68", -- 0x1B38
    x"F0",x"20",x"C9",x"64",x"F0",x"03",x"20",x"77", -- 0x1B40
    x"DA",x"84",x"99",x"68",x"4A",x"85",x"63",x"68", -- 0x1B48
    x"85",x"B3",x"68",x"85",x"B4",x"68",x"85",x"B5", -- 0x1B50
    x"68",x"85",x"B6",x"68",x"85",x"B7",x"45",x"B0", -- 0x1B58
    x"85",x"B8",x"A5",x"AC",x"60",x"A5",x"C3",x"A4", -- 0x1B60
    x"C4",x"69",x"00",x"90",x"01",x"C8",x"20",x"EB", -- 0x1B68
    x"E0",x"4C",x"76",x"E4",x"20",x"BC",x"00",x"B0", -- 0x1B70
    x"03",x"4C",x"50",x"E9",x"AA",x"30",x"2F",x"C9", -- 0x1B78
    x"24",x"F0",x"F6",x"C9",x"25",x"F0",x"F2",x"C9", -- 0x1B80
    x"2E",x"F0",x"EE",x"C9",x"22",x"F0",x"D6",x"C9", -- 0x1B88
    x"28",x"D0",x"4F",x"20",x"90",x"DA",x"A9",x"29", -- 0x1B90
    x"A0",x"00",x"D1",x"C3",x"D0",x"0B",x"4C",x"BC", -- 0x1B98
    x"00",x"A9",x"28",x"D0",x"F3",x"A9",x"2C",x"D0", -- 0x1BA0
    x"EF",x"A2",x"02",x"4C",x"2B",x"D1",x"C9",x"B6", -- 0x1BA8
    x"F0",x"29",x"C9",x"B5",x"F0",x"BE",x"C9",x"B0", -- 0x1BB0
    x"D0",x"13",x"A0",x"21",x"D0",x"1F",x"20",x"4D", -- 0x1BB8
    x"DE",x"A5",x"AF",x"49",x"FF",x"A8",x"A5",x"AE", -- 0x1BC0
    x"49",x"FF",x"4C",x"00",x"E0",x"C9",x"AD",x"D0", -- 0x1BC8
    x"03",x"4C",x"5B",x"E0",x"E9",x"C2",x"B0",x"19", -- 0x1BD0
    x"4C",x"A9",x"DB",x"A0",x"1E",x"68",x"68",x"4C", -- 0x1BD8
    x"E1",x"DA",x"20",x"51",x"DD",x"85",x"AE",x"84", -- 0x1BE0
    x"AF",x"A6",x"5F",x"30",x"03",x"4C",x"27",x"E8", -- 0x1BE8
    x"60",x"0A",x"A8",x"B9",x"4A",x"F2",x"48",x"B9", -- 0x1BF0
    x"49",x"F2",x"48",x"B9",x"04",x"F2",x"F0",x"05", -- 0x1BF8
    x"48",x"B9",x"03",x"F2",x"48",x"60",x"20",x"93", -- 0x1C00
    x"DB",x"4C",x"79",x"DA",x"20",x"93",x"DB",x"4C", -- 0x1C08
    x"77",x"DA",x"46",x"5F",x"4C",x"BC",x"00",x"20", -- 0x1C10
    x"90",x"DA",x"20",x"A5",x"DB",x"20",x"79",x"DA", -- 0x1C18
    x"68",x"AA",x"68",x"A8",x"A5",x"AF",x"48",x"A5", -- 0x1C20
    x"AE",x"48",x"98",x"48",x"8A",x"48",x"20",x"33", -- 0x1C28
    x"E4",x"8A",x"60",x"20",x"90",x"DA",x"20",x"77", -- 0x1C30
    x"DA",x"A5",x"AC",x"C9",x"98",x"B0",x"20",x"20", -- 0x1C38
    x"FA",x"E8",x"A2",x"02",x"B5",x"AD",x"95",x"11", -- 0x1C40
    x"CA",x"10",x"F9",x"20",x"C2",x"00",x"A2",x"00", -- 0x1C48
    x"C9",x"29",x"F0",x"0A",x"20",x"85",x"E4",x"20", -- 0x1C50
    x"C2",x"00",x"C9",x"29",x"D0",x"01",x"60",x"4C", -- 0x1C58
    x"D0",x"DE",x"20",x"89",x"DC",x"45",x"5B",x"A8", -- 0x1C60
    x"A5",x"AE",x"45",x"5C",x"4C",x"00",x"E0",x"20", -- 0x1C68
    x"89",x"DC",x"05",x"5B",x"A8",x"A5",x"AE",x"05", -- 0x1C70
    x"5C",x"4C",x"00",x"E0",x"20",x"89",x"DC",x"25", -- 0x1C78
    x"5B",x"A8",x"A5",x"AE",x"25",x"5C",x"4C",x"00", -- 0x1C80
    x"E0",x"20",x"4D",x"DE",x"A5",x"AE",x"85",x"5C", -- 0x1C88
    x"A5",x"AF",x"85",x"5B",x"20",x"6A",x"E5",x"20", -- 0x1C90
    x"4D",x"DE",x"A5",x"AF",x"60",x"20",x"7A",x"DA", -- 0x1C98
    x"B0",x"13",x"A5",x"B7",x"09",x"7F",x"25",x"B4", -- 0x1CA0
    x"85",x"B4",x"A9",x"B3",x"A0",x"00",x"20",x"C1", -- 0x1CA8
    x"E8",x"AA",x"4C",x"E6",x"DC",x"46",x"5F",x"C6", -- 0x1CB0
    x"9B",x"20",x"E5",x"E2",x"85",x"AC",x"86",x"AD", -- 0x1CB8
    x"84",x"AE",x"A5",x"B5",x"A4",x"B6",x"20",x"E9", -- 0x1CC0
    x"E2",x"86",x"B5",x"84",x"B6",x"AA",x"38",x"E5", -- 0x1CC8
    x"AC",x"F0",x"08",x"A9",x"01",x"90",x"04",x"A6", -- 0x1CD0
    x"AC",x"A9",x"FF",x"85",x"B0",x"A0",x"FF",x"E8", -- 0x1CD8
    x"C8",x"CA",x"D0",x"07",x"A6",x"B0",x"30",x"0F", -- 0x1CE0
    x"18",x"90",x"0C",x"B1",x"B5",x"D1",x"AD",x"F0", -- 0x1CE8
    x"EF",x"A2",x"FF",x"B0",x"02",x"A2",x"01",x"E8", -- 0x1CF0
    x"8A",x"2A",x"25",x"63",x"F0",x"02",x"A9",x"FF", -- 0x1CF8
    x"4C",x"A4",x"E8",x"20",x"A5",x"DB",x"AA",x"20", -- 0x1D00
    x"56",x"DD",x"20",x"C2",x"00",x"D0",x"F4",x"60", -- 0x1D08
    x"20",x"46",x"DD",x"A5",x"AE",x"A6",x"78",x"F0", -- 0x1D10
    x"22",x"E0",x"10",x"B0",x"23",x"06",x"AF",x"2A", -- 0x1D18
    x"CA",x"D0",x"FA",x"A4",x"AF",x"4C",x"00",x"E0", -- 0x1D20
    x"20",x"46",x"DD",x"A5",x"AE",x"A6",x"78",x"F0", -- 0x1D28
    x"0A",x"E0",x"10",x"B0",x"0B",x"4A",x"66",x"AF", -- 0x1D30
    x"CA",x"D0",x"FA",x"A4",x"AF",x"4C",x"00",x"E0", -- 0x1D38
    x"A9",x"00",x"A8",x"4C",x"00",x"E0",x"20",x"36", -- 0x1D40
    x"E4",x"86",x"78",x"20",x"6A",x"E5",x"4C",x"4D", -- 0x1D48
    x"DE",x"A2",x"00",x"20",x"C2",x"00",x"86",x"5E", -- 0x1D50
    x"85",x"93",x"29",x"7F",x"20",x"C5",x"DD",x"B0", -- 0x1D58
    x"03",x"4C",x"A9",x"DB",x"A2",x"00",x"86",x"5F", -- 0x1D60
    x"20",x"BC",x"00",x"90",x"05",x"20",x"C5",x"DD", -- 0x1D68
    x"90",x"0B",x"AA",x"20",x"BC",x"00",x"90",x"FB", -- 0x1D70
    x"20",x"C5",x"DD",x"B0",x"F6",x"C9",x"24",x"D0", -- 0x1D78
    x"0B",x"A9",x"FF",x"85",x"5F",x"8A",x"09",x"80", -- 0x1D80
    x"AA",x"20",x"BC",x"00",x"86",x"94",x"05",x"61", -- 0x1D88
    x"C9",x"28",x"D0",x"03",x"4C",x"5F",x"DE",x"A9", -- 0x1D90
    x"00",x"85",x"61",x"A5",x"7B",x"A6",x"7C",x"A0", -- 0x1D98
    x"00",x"86",x"AB",x"85",x"AA",x"E4",x"7E",x"D0", -- 0x1DA0
    x"04",x"C5",x"7D",x"F0",x"2C",x"A5",x"93",x"D1", -- 0x1DA8
    x"AA",x"D0",x"08",x"A5",x"94",x"C8",x"D1",x"AA", -- 0x1DB0
    x"F0",x"69",x"88",x"18",x"A5",x"AA",x"69",x"06", -- 0x1DB8
    x"90",x"E1",x"E8",x"D0",x"DC",x"C9",x"61",x"B0", -- 0x1DC0
    x"0A",x"C9",x"41",x"90",x"05",x"E9",x"5B",x"38", -- 0x1DC8
    x"E9",x"A5",x"60",x"E9",x"7B",x"38",x"E9",x"85", -- 0x1DD0
    x"60",x"68",x"48",x"C9",x"E4",x"D0",x"05",x"A9", -- 0x1DD8
    x"87",x"A0",x"F1",x"60",x"A5",x"7D",x"A4",x"7E", -- 0x1DE0
    x"85",x"AA",x"84",x"AB",x"A5",x"7F",x"A4",x"80", -- 0x1DE8
    x"85",x"A6",x"84",x"A7",x"18",x"69",x"06",x"90", -- 0x1DF0
    x"01",x"C8",x"85",x"A4",x"84",x"A5",x"20",x"B2", -- 0x1DF8
    x"D0",x"A5",x"A4",x"A4",x"A5",x"C8",x"85",x"7D", -- 0x1E00
    x"84",x"7E",x"A0",x"00",x"A5",x"93",x"91",x"AA", -- 0x1E08
    x"C8",x"A5",x"94",x"91",x"AA",x"A9",x"00",x"C8", -- 0x1E10
    x"91",x"AA",x"C8",x"91",x"AA",x"C8",x"91",x"AA", -- 0x1E18
    x"C8",x"91",x"AA",x"A5",x"AA",x"18",x"69",x"02", -- 0x1E20
    x"A4",x"AB",x"90",x"01",x"C8",x"85",x"95",x"84", -- 0x1E28
    x"96",x"60",x"A5",x"5D",x"0A",x"69",x"05",x"65", -- 0x1E30
    x"AA",x"A4",x"AB",x"90",x"01",x"C8",x"85",x"A4", -- 0x1E38
    x"84",x"A5",x"60",x"20",x"BC",x"00",x"20",x"74", -- 0x1E40
    x"DA",x"A5",x"B0",x"30",x"0D",x"A5",x"AC",x"C9", -- 0x1E48
    x"90",x"90",x"09",x"A9",x"8E",x"A0",x"F1",x"20", -- 0x1E50
    x"C1",x"E8",x"D0",x"74",x"4C",x"FA",x"E8",x"A5", -- 0x1E58
    x"5E",x"48",x"A5",x"5F",x"48",x"A0",x"00",x"98", -- 0x1E60
    x"48",x"A5",x"94",x"48",x"A5",x"93",x"48",x"20", -- 0x1E68
    x"43",x"DE",x"68",x"85",x"93",x"68",x"85",x"94", -- 0x1E70
    x"68",x"A8",x"BA",x"BD",x"02",x"01",x"48",x"BD", -- 0x1E78
    x"01",x"01",x"48",x"A5",x"AE",x"9D",x"02",x"01", -- 0x1E80
    x"A5",x"AF",x"9D",x"01",x"01",x"C8",x"20",x"C2", -- 0x1E88
    x"00",x"C9",x"2C",x"F0",x"D2",x"84",x"5D",x"20", -- 0x1E90
    x"96",x"DB",x"68",x"85",x"5F",x"68",x"85",x"5E", -- 0x1E98
    x"A6",x"7D",x"A5",x"7E",x"86",x"AA",x"85",x"AB", -- 0x1EA0
    x"C5",x"80",x"D0",x"04",x"E4",x"7F",x"F0",x"39", -- 0x1EA8
    x"A0",x"00",x"B1",x"AA",x"C8",x"C5",x"93",x"D0", -- 0x1EB0
    x"06",x"A5",x"94",x"D1",x"AA",x"F0",x"16",x"C8", -- 0x1EB8
    x"B1",x"AA",x"18",x"65",x"AA",x"AA",x"C8",x"B1", -- 0x1EC0
    x"AA",x"65",x"AB",x"90",x"D7",x"A2",x"10",x"2C", -- 0x1EC8
    x"A2",x"08",x"4C",x"2B",x"D1",x"A2",x"12",x"A5", -- 0x1ED0
    x"5E",x"D0",x"F7",x"20",x"32",x"DE",x"A5",x"5D", -- 0x1ED8
    x"A0",x"04",x"D1",x"AA",x"D0",x"E7",x"4C",x"6C", -- 0x1EE0
    x"DF",x"20",x"32",x"DE",x"20",x"FC",x"D0",x"A0", -- 0x1EE8
    x"00",x"84",x"BB",x"A5",x"93",x"91",x"AA",x"C8", -- 0x1EF0
    x"A5",x"94",x"91",x"AA",x"A5",x"5D",x"A0",x"04", -- 0x1EF8
    x"84",x"BA",x"91",x"AA",x"18",x"A2",x"0B",x"A9", -- 0x1F00
    x"00",x"24",x"5E",x"50",x"07",x"68",x"69",x"01", -- 0x1F08
    x"AA",x"68",x"69",x"00",x"C8",x"91",x"AA",x"C8", -- 0x1F10
    x"8A",x"91",x"AA",x"20",x"BB",x"DF",x"86",x"BA", -- 0x1F18
    x"85",x"BB",x"A4",x"71",x"C6",x"5D",x"D0",x"DD", -- 0x1F20
    x"65",x"A5",x"B0",x"5D",x"85",x"A5",x"A8",x"8A", -- 0x1F28
    x"65",x"A4",x"90",x"03",x"C8",x"F0",x"52",x"20", -- 0x1F30
    x"FC",x"D0",x"85",x"7F",x"84",x"80",x"A9",x"00", -- 0x1F38
    x"E6",x"BB",x"A4",x"BA",x"F0",x"05",x"88",x"91", -- 0x1F40
    x"A4",x"D0",x"FB",x"C6",x"A5",x"C6",x"BB",x"D0", -- 0x1F48
    x"F5",x"E6",x"A5",x"38",x"A0",x"02",x"A5",x"7F", -- 0x1F50
    x"E5",x"AA",x"91",x"AA",x"C8",x"A5",x"80",x"E5", -- 0x1F58
    x"AB",x"91",x"AA",x"A5",x"5E",x"D0",x"53",x"C8", -- 0x1F60
    x"B1",x"AA",x"85",x"5D",x"A9",x"00",x"85",x"BA", -- 0x1F68
    x"85",x"BB",x"C8",x"68",x"AA",x"85",x"AE",x"68", -- 0x1F70
    x"85",x"AF",x"D1",x"AA",x"90",x"0E",x"D0",x"06", -- 0x1F78
    x"C8",x"8A",x"D1",x"AA",x"90",x"07",x"4C",x"CD", -- 0x1F80
    x"DE",x"4C",x"29",x"D1",x"C8",x"A5",x"BB",x"05", -- 0x1F88
    x"BA",x"F0",x"0A",x"20",x"BB",x"DF",x"8A",x"65", -- 0x1F90
    x"AE",x"AA",x"98",x"A4",x"71",x"65",x"AF",x"86", -- 0x1F98
    x"BA",x"C6",x"5D",x"D0",x"CB",x"06",x"BA",x"2A", -- 0x1FA0
    x"06",x"BA",x"2A",x"A8",x"A5",x"BA",x"65",x"A4", -- 0x1FA8
    x"85",x"95",x"98",x"65",x"A5",x"85",x"96",x"A8", -- 0x1FB0
    x"A5",x"95",x"60",x"84",x"71",x"B1",x"AA",x"85", -- 0x1FB8
    x"76",x"88",x"B1",x"AA",x"85",x"77",x"A9",x"10", -- 0x1FC0
    x"85",x"A8",x"A2",x"00",x"A0",x"00",x"8A",x"0A", -- 0x1FC8
    x"AA",x"98",x"2A",x"A8",x"B0",x"B3",x"06",x"BA", -- 0x1FD0
    x"26",x"BB",x"90",x"0B",x"18",x"8A",x"65",x"76", -- 0x1FD8
    x"AA",x"98",x"65",x"77",x"A8",x"B0",x"A2",x"C6", -- 0x1FE0
    x"A8",x"D0",x"E3",x"60",x"A5",x"5F",x"10",x"03", -- 0x1FE8
    x"20",x"E5",x"E2",x"20",x"86",x"E1",x"38",x"A5", -- 0x1FF0
    x"81",x"E5",x"7F",x"A8",x"A5",x"82",x"E5",x"80", -- 0x1FF8
    x"46",x"5F",x"85",x"AD",x"84",x"AE",x"A2",x"90", -- 0x2000
    x"4C",x"AC",x"E8",x"A4",x"0E",x"A9",x"00",x"F0", -- 0x2008
    x"EF",x"A6",x"88",x"E8",x"D0",x"A4",x"A2",x"16", -- 0x2010
    x"4C",x"2B",x"D1",x"20",x"4C",x"E0",x"85",x"9C", -- 0x2018
    x"84",x"9D",x"20",x"11",x"E0",x"20",x"A1",x"DB", -- 0x2020
    x"A9",x"80",x"85",x"61",x"20",x"51",x"DD",x"20", -- 0x2028
    x"77",x"DA",x"20",x"96",x"DB",x"A9",x"C0",x"20", -- 0x2030
    x"98",x"DB",x"A5",x"96",x"48",x"A5",x"95",x"48", -- 0x2038
    x"A5",x"C4",x"48",x"A5",x"C3",x"48",x"20",x"7B", -- 0x2040
    x"D6",x"4C",x"BB",x"E0",x"A9",x"AD",x"20",x"98", -- 0x2048
    x"DB",x"09",x"80",x"85",x"61",x"20",x"58",x"DD", -- 0x2050
    x"4C",x"77",x"DA",x"20",x"4C",x"E0",x"48",x"98", -- 0x2058
    x"48",x"20",x"A1",x"DB",x"20",x"88",x"DA",x"20", -- 0x2060
    x"96",x"DB",x"20",x"77",x"DA",x"68",x"85",x"9D", -- 0x2068
    x"68",x"85",x"9C",x"A2",x"20",x"A0",x"03",x"B1", -- 0x2070
    x"9C",x"F0",x"9D",x"85",x"96",x"88",x"B1",x"9C", -- 0x2078
    x"85",x"95",x"AA",x"C8",x"B1",x"95",x"48",x"88", -- 0x2080
    x"10",x"FA",x"A4",x"96",x"20",x"51",x"E8",x"A5", -- 0x2088
    x"C4",x"48",x"A5",x"C3",x"48",x"B1",x"9C",x"85", -- 0x2090
    x"C3",x"C8",x"B1",x"9C",x"85",x"C4",x"A5",x"96", -- 0x2098
    x"48",x"A5",x"95",x"48",x"20",x"74",x"DA",x"68", -- 0x20A0
    x"85",x"9C",x"68",x"85",x"9D",x"20",x"C2",x"00", -- 0x20A8
    x"F0",x"03",x"4C",x"A9",x"DB",x"68",x"85",x"C3", -- 0x20B0
    x"68",x"85",x"C4",x"A0",x"00",x"68",x"91",x"9C", -- 0x20B8
    x"C8",x"68",x"91",x"9C",x"C8",x"68",x"91",x"9C", -- 0x20C0
    x"C8",x"68",x"91",x"9C",x"60",x"20",x"77",x"DA", -- 0x20C8
    x"20",x"40",x"EA",x"A9",x"F0",x"A0",x"00",x"F0", -- 0x20D0
    x"12",x"A6",x"AE",x"A4",x"AF",x"86",x"9E",x"84", -- 0x20D8
    x"9F",x"20",x"54",x"E1",x"86",x"AD",x"84",x"AE", -- 0x20E0
    x"85",x"AC",x"60",x"A2",x"22",x"86",x"5B",x"86", -- 0x20E8
    x"5C",x"85",x"B8",x"84",x"B9",x"85",x"AD",x"84", -- 0x20F0
    x"AE",x"A0",x"FF",x"C8",x"B1",x"B8",x"F0",x"0C", -- 0x20F8
    x"C5",x"5B",x"F0",x"04",x"C5",x"5C",x"D0",x"F3", -- 0x2100
    x"C9",x"22",x"F0",x"01",x"18",x"84",x"AC",x"98", -- 0x2108
    x"65",x"B8",x"85",x"BA",x"A6",x"B9",x"90",x"01", -- 0x2110
    x"E8",x"86",x"BB",x"A5",x"B9",x"C9",x"04",x"B0", -- 0x2118
    x"0B",x"98",x"20",x"D9",x"E0",x"A6",x"B8",x"A4", -- 0x2120
    x"B9",x"20",x"C6",x"E2",x"A6",x"65",x"E0",x"71", -- 0x2128
    x"D0",x"05",x"A2",x"1C",x"4C",x"2B",x"D1",x"A5", -- 0x2130
    x"AC",x"95",x"00",x"A5",x"AD",x"95",x"01",x"A5", -- 0x2138
    x"AE",x"95",x"02",x"A0",x"00",x"86",x"AE",x"84", -- 0x2140
    x"AF",x"88",x"84",x"5F",x"86",x"66",x"E8",x"E8", -- 0x2148
    x"E8",x"86",x"65",x"60",x"46",x"60",x"48",x"49", -- 0x2150
    x"FF",x"38",x"65",x"81",x"A4",x"82",x"B0",x"01", -- 0x2158
    x"88",x"C4",x"80",x"90",x"11",x"D0",x"04",x"C5", -- 0x2160
    x"7F",x"90",x"0B",x"85",x"81",x"84",x"82",x"85", -- 0x2168
    x"83",x"84",x"84",x"AA",x"68",x"60",x"A2",x"0C", -- 0x2170
    x"A5",x"60",x"30",x"B8",x"20",x"86",x"E1",x"A9", -- 0x2178
    x"80",x"85",x"60",x"68",x"D0",x"D0",x"A6",x"85", -- 0x2180
    x"A5",x"86",x"86",x"81",x"85",x"82",x"A0",x"00", -- 0x2188
    x"84",x"9D",x"A5",x"7F",x"A6",x"80",x"85",x"AA", -- 0x2190
    x"86",x"AB",x"A9",x"68",x"85",x"71",x"84",x"72", -- 0x2198
    x"C5",x"65",x"F0",x"05",x"20",x"0A",x"E2",x"F0", -- 0x21A0
    x"F7",x"06",x"A0",x"A5",x"7B",x"A6",x"7C",x"85", -- 0x21A8
    x"71",x"86",x"72",x"E4",x"7E",x"D0",x"04",x"C5", -- 0x21B0
    x"7D",x"F0",x"05",x"20",x"04",x"E2",x"F0",x"F3", -- 0x21B8
    x"85",x"A4",x"86",x"A5",x"A9",x"04",x"85",x"A0", -- 0x21C0
    x"A5",x"A4",x"A6",x"A5",x"E4",x"80",x"D0",x"04", -- 0x21C8
    x"C5",x"7F",x"F0",x"75",x"85",x"71",x"86",x"72", -- 0x21D0
    x"A0",x"02",x"B1",x"71",x"65",x"A4",x"85",x"A4", -- 0x21D8
    x"C8",x"B1",x"71",x"65",x"A5",x"85",x"A5",x"A0", -- 0x21E0
    x"01",x"B1",x"71",x"10",x"DB",x"A0",x"04",x"B1", -- 0x21E8
    x"71",x"0A",x"69",x"05",x"20",x"3C",x"E2",x"E4", -- 0x21F0
    x"A5",x"D0",x"04",x"C5",x"A4",x"F0",x"CD",x"20", -- 0x21F8
    x"0A",x"E2",x"F0",x"F3",x"C8",x"B1",x"71",x"10", -- 0x2200
    x"30",x"C8",x"B1",x"71",x"F0",x"2B",x"C8",x"B1", -- 0x2208
    x"71",x"AA",x"C8",x"B1",x"71",x"C5",x"82",x"90", -- 0x2210
    x"06",x"D0",x"1E",x"E4",x"81",x"B0",x"1A",x"C5", -- 0x2218
    x"AB",x"90",x"17",x"D0",x"04",x"E4",x"AA",x"90", -- 0x2220
    x"11",x"86",x"AA",x"85",x"AB",x"A5",x"71",x"A6", -- 0x2228
    x"72",x"85",x"9C",x"86",x"9D",x"88",x"88",x"84", -- 0x2230
    x"A2",x"18",x"A5",x"A0",x"65",x"71",x"85",x"71", -- 0x2238
    x"90",x"02",x"E6",x"72",x"A6",x"72",x"A0",x"00", -- 0x2240
    x"60",x"C6",x"A0",x"A6",x"9D",x"F0",x"F5",x"A4", -- 0x2248
    x"A2",x"18",x"B1",x"9C",x"65",x"AA",x"85",x"A6", -- 0x2250
    x"A5",x"AB",x"69",x"00",x"85",x"A7",x"A5",x"81", -- 0x2258
    x"A6",x"82",x"85",x"A4",x"86",x"A5",x"20",x"B9", -- 0x2260
    x"D0",x"A4",x"A2",x"C8",x"A5",x"A4",x"91",x"9C", -- 0x2268
    x"AA",x"E6",x"A5",x"A5",x"A5",x"C8",x"91",x"9C", -- 0x2270
    x"4C",x"8A",x"E1",x"A5",x"AF",x"48",x"A5",x"AE", -- 0x2278
    x"48",x"20",x"74",x"DB",x"20",x"79",x"DA",x"68", -- 0x2280
    x"85",x"B8",x"68",x"85",x"B9",x"A0",x"00",x"B1", -- 0x2288
    x"B8",x"18",x"71",x"AE",x"90",x"05",x"A2",x"1A", -- 0x2290
    x"4C",x"2B",x"D1",x"20",x"D9",x"E0",x"20",x"B8", -- 0x2298
    x"E2",x"A5",x"9E",x"A4",x"9F",x"20",x"E9",x"E2", -- 0x22A0
    x"20",x"CA",x"E2",x"A5",x"B8",x"A4",x"B9",x"20", -- 0x22A8
    x"E9",x"E2",x"20",x"2C",x"E1",x"4C",x"9F",x"DA", -- 0x22B0
    x"A0",x"00",x"B1",x"B8",x"48",x"C8",x"B1",x"B8", -- 0x22B8
    x"AA",x"C8",x"B1",x"B8",x"A8",x"68",x"86",x"71", -- 0x22C0
    x"84",x"72",x"AA",x"F0",x"14",x"A0",x"00",x"B1", -- 0x22C8
    x"71",x"91",x"83",x"C8",x"CA",x"D0",x"F8",x"98", -- 0x22D0
    x"18",x"65",x"83",x"85",x"83",x"90",x"02",x"E6", -- 0x22D8
    x"84",x"60",x"20",x"79",x"DA",x"A5",x"AE",x"A4", -- 0x22E0
    x"AF",x"85",x"71",x"84",x"72",x"20",x"1A",x"E3", -- 0x22E8
    x"08",x"A0",x"00",x"B1",x"71",x"48",x"C8",x"B1", -- 0x22F0
    x"71",x"AA",x"C8",x"B1",x"71",x"A8",x"68",x"28", -- 0x22F8
    x"D0",x"13",x"C4",x"82",x"D0",x"0F",x"E4",x"81", -- 0x2300
    x"D0",x"0B",x"48",x"18",x"65",x"81",x"85",x"81", -- 0x2308
    x"90",x"02",x"E6",x"82",x"68",x"86",x"71",x"84", -- 0x2310
    x"72",x"60",x"C4",x"67",x"D0",x"0C",x"C5",x"66", -- 0x2318
    x"D0",x"08",x"85",x"65",x"E9",x"03",x"85",x"66", -- 0x2320
    x"A0",x"00",x"60",x"20",x"36",x"E4",x"8A",x"48", -- 0x2328
    x"A9",x"01",x"20",x"E1",x"E0",x"68",x"A0",x"00", -- 0x2330
    x"91",x"AD",x"4C",x"2C",x"E1",x"48",x"20",x"9E", -- 0x2338
    x"E3",x"D1",x"9E",x"98",x"F0",x"09",x"48",x"20", -- 0x2340
    x"9E",x"E3",x"18",x"F1",x"9E",x"49",x"FF",x"90", -- 0x2348
    x"04",x"B1",x"9E",x"AA",x"98",x"48",x"8A",x"48", -- 0x2350
    x"20",x"E1",x"E0",x"A5",x"9E",x"A4",x"9F",x"20", -- 0x2358
    x"E9",x"E2",x"68",x"A8",x"68",x"18",x"65",x"71", -- 0x2360
    x"85",x"71",x"90",x"02",x"E6",x"72",x"98",x"20", -- 0x2368
    x"CA",x"E2",x"4C",x"2C",x"E1",x"48",x"A9",x"FF", -- 0x2370
    x"85",x"AF",x"20",x"C2",x"00",x"C9",x"29",x"F0", -- 0x2378
    x"06",x"20",x"A5",x"DB",x"20",x"33",x"E4",x"20", -- 0x2380
    x"9E",x"E3",x"CA",x"8A",x"48",x"18",x"A2",x"00", -- 0x2388
    x"F1",x"9E",x"B0",x"C2",x"49",x"FF",x"C5",x"AF", -- 0x2390
    x"90",x"BD",x"A5",x"AF",x"B0",x"B9",x"20",x"96", -- 0x2398
    x"DB",x"68",x"85",x"A2",x"68",x"85",x"A3",x"68", -- 0x23A0
    x"AA",x"68",x"85",x"9E",x"68",x"85",x"9F",x"A0", -- 0x23A8
    x"00",x"8A",x"F0",x"79",x"E6",x"A2",x"6C",x"A2", -- 0x23B0
    x"00",x"20",x"E2",x"E2",x"85",x"AC",x"A8",x"F0", -- 0x23B8
    x"38",x"20",x"E1",x"E0",x"86",x"AD",x"84",x"AE", -- 0x23C0
    x"A8",x"88",x"B1",x"71",x"20",x"C9",x"DD",x"90", -- 0x23C8
    x"02",x"09",x"20",x"91",x"83",x"98",x"D0",x"F1", -- 0x23D0
    x"F0",x"1F",x"20",x"E2",x"E2",x"85",x"AC",x"A8", -- 0x23D8
    x"F0",x"17",x"20",x"E1",x"E0",x"86",x"AD",x"84", -- 0x23E0
    x"AE",x"A8",x"88",x"B1",x"71",x"20",x"C5",x"DD", -- 0x23E8
    x"90",x"02",x"29",x"DF",x"91",x"83",x"98",x"D0", -- 0x23F0
    x"F1",x"4C",x"2C",x"E1",x"20",x"BC",x"00",x"20", -- 0x23F8
    x"51",x"DD",x"20",x"96",x"DB",x"20",x"79",x"DA", -- 0x2400
    x"A0",x"02",x"B1",x"95",x"AA",x"88",x"B1",x"95", -- 0x2408
    x"A8",x"8A",x"4C",x"00",x"E0",x"20",x"1B",x"E4", -- 0x2410
    x"4C",x"0D",x"E0",x"20",x"E2",x"E2",x"A8",x"60", -- 0x2418
    x"20",x"1B",x"E4",x"F0",x"08",x"A0",x"00",x"B1", -- 0x2420
    x"71",x"A8",x"4C",x"0D",x"E0",x"4C",x"D0",x"DE", -- 0x2428
    x"20",x"BC",x"00",x"20",x"74",x"DA",x"20",x"49", -- 0x2430
    x"DE",x"A4",x"AE",x"D0",x"F0",x"A6",x"AF",x"4C", -- 0x2438
    x"C2",x"00",x"20",x"1B",x"E4",x"D0",x"03",x"4C", -- 0x2440
    x"F7",x"E5",x"A6",x"C3",x"A4",x"C4",x"86",x"BA", -- 0x2448
    x"84",x"BB",x"A6",x"71",x"86",x"C3",x"18",x"65", -- 0x2450
    x"71",x"85",x"73",x"A5",x"72",x"85",x"C4",x"69", -- 0x2458
    x"00",x"85",x"74",x"A0",x"00",x"B1",x"73",x"48", -- 0x2460
    x"98",x"91",x"73",x"20",x"C2",x"00",x"20",x"50", -- 0x2468
    x"E9",x"68",x"A0",x"00",x"91",x"73",x"A6",x"BA", -- 0x2470
    x"A4",x"BB",x"86",x"C3",x"84",x"C4",x"60",x"20", -- 0x2478
    x"74",x"DA",x"20",x"98",x"E4",x"20",x"A5",x"DB", -- 0x2480
    x"A5",x"12",x"48",x"A5",x"11",x"48",x"20",x"33", -- 0x2488
    x"E4",x"68",x"85",x"11",x"68",x"85",x"12",x"60", -- 0x2490
    x"A5",x"AC",x"C9",x"98",x"B0",x"8F",x"20",x"FA", -- 0x2498
    x"E8",x"A5",x"AE",x"A4",x"AF",x"84",x"11",x"85", -- 0x24A0
    x"12",x"60",x"20",x"98",x"E4",x"A2",x"00",x"A1", -- 0x24A8
    x"11",x"A8",x"4C",x"0D",x"E0",x"20",x"7F",x"E4", -- 0x24B0
    x"8A",x"A2",x"00",x"81",x"11",x"60",x"20",x"98", -- 0x24B8
    x"E4",x"A2",x"00",x"A1",x"11",x"A8",x"E6",x"11", -- 0x24C0
    x"D0",x"02",x"E6",x"12",x"A1",x"11",x"4C",x"00", -- 0x24C8
    x"E0",x"20",x"74",x"DA",x"20",x"98",x"E4",x"84", -- 0x24D0
    x"97",x"85",x"98",x"20",x"A5",x"DB",x"20",x"74", -- 0x24D8
    x"DA",x"20",x"98",x"E4",x"98",x"A2",x"00",x"81", -- 0x24E0
    x"97",x"E6",x"97",x"D0",x"02",x"E6",x"98",x"A5", -- 0x24E8
    x"12",x"81",x"97",x"4C",x"C2",x"00",x"20",x"51", -- 0x24F0
    x"DD",x"85",x"97",x"84",x"98",x"A5",x"5F",x"48", -- 0x24F8
    x"20",x"A5",x"DB",x"20",x"51",x"DD",x"68",x"45", -- 0x2500
    x"5F",x"10",x"10",x"A0",x"03",x"B1",x"97",x"48", -- 0x2508
    x"B1",x"95",x"91",x"97",x"68",x"91",x"95",x"88", -- 0x2510
    x"10",x"F3",x"60",x"4C",x"83",x"DA",x"20",x"74", -- 0x2518
    x"DA",x"20",x"98",x"E4",x"A9",x"E5",x"48",x"A9", -- 0x2520
    x"2C",x"48",x"6C",x"11",x"00",x"4C",x"C2",x"00", -- 0x2528
    x"20",x"7F",x"E4",x"86",x"97",x"A2",x"00",x"20", -- 0x2530
    x"C2",x"00",x"F0",x"03",x"20",x"85",x"E4",x"86", -- 0x2538
    x"98",x"B1",x"11",x"45",x"98",x"25",x"97",x"F0", -- 0x2540
    x"F8",x"60",x"20",x"32",x"E7",x"A5",x"B0",x"49", -- 0x2548
    x"FF",x"85",x"B0",x"45",x"B7",x"85",x"B8",x"A5", -- 0x2550
    x"AC",x"4C",x"68",x"E5",x"20",x"81",x"E6",x"90", -- 0x2558
    x"4D",x"A9",x"8F",x"A0",x"F1",x"20",x"32",x"E7", -- 0x2560
    x"D0",x"10",x"A5",x"B7",x"85",x"B0",x"A2",x"04", -- 0x2568
    x"B5",x"B2",x"95",x"AB",x"CA",x"D0",x"F9",x"86", -- 0x2570
    x"B9",x"60",x"A6",x"B9",x"86",x"A3",x"A2",x"B3", -- 0x2578
    x"A5",x"B3",x"A8",x"F0",x"C4",x"38",x"E5",x"AC", -- 0x2580
    x"F0",x"24",x"90",x"12",x"84",x"AC",x"A4",x"B7", -- 0x2588
    x"84",x"B0",x"49",x"FF",x"69",x"00",x"A0",x"00", -- 0x2590
    x"84",x"A3",x"A2",x"AC",x"D0",x"04",x"A0",x"00", -- 0x2598
    x"84",x"B9",x"C9",x"F9",x"30",x"B6",x"A8",x"A5", -- 0x25A0
    x"B9",x"56",x"01",x"20",x"98",x"E6",x"24",x"B8", -- 0x25A8
    x"10",x"4C",x"A0",x"AC",x"E0",x"B3",x"F0",x"02", -- 0x25B0
    x"A0",x"B3",x"38",x"49",x"FF",x"65",x"A3",x"85", -- 0x25B8
    x"B9",x"B9",x"03",x"00",x"F5",x"03",x"85",x"AF", -- 0x25C0
    x"B9",x"02",x"00",x"F5",x"02",x"85",x"AE",x"B9", -- 0x25C8
    x"01",x"00",x"F5",x"01",x"85",x"AD",x"B0",x"03", -- 0x25D0
    x"20",x"3D",x"E6",x"A0",x"00",x"98",x"18",x"A6", -- 0x25D8
    x"AD",x"D0",x"3E",x"A6",x"AE",x"86",x"AD",x"A6", -- 0x25E0
    x"AF",x"86",x"AE",x"A6",x"B9",x"86",x"AF",x"84", -- 0x25E8
    x"B9",x"69",x"08",x"C9",x"18",x"D0",x"E8",x"A9", -- 0x25F0
    x"00",x"85",x"AC",x"85",x"B0",x"60",x"65",x"A3", -- 0x25F8
    x"85",x"B9",x"A5",x"AF",x"65",x"B6",x"85",x"AF", -- 0x2600
    x"A5",x"AE",x"65",x"B5",x"85",x"AE",x"A5",x"AD", -- 0x2608
    x"65",x"B4",x"85",x"AD",x"B0",x"1A",x"60",x"69", -- 0x2610
    x"01",x"06",x"B9",x"26",x"AF",x"26",x"AE",x"26", -- 0x2618
    x"AD",x"10",x"F4",x"38",x"E5",x"AC",x"B0",x"CF", -- 0x2620
    x"49",x"FF",x"69",x"01",x"85",x"AC",x"90",x"0C", -- 0x2628
    x"E6",x"AC",x"F0",x"36",x"66",x"AD",x"66",x"AE", -- 0x2630
    x"66",x"AF",x"66",x"B9",x"60",x"A5",x"B0",x"49", -- 0x2638
    x"FF",x"85",x"B0",x"A5",x"AD",x"49",x"FF",x"85", -- 0x2640
    x"AD",x"A5",x"AE",x"49",x"FF",x"85",x"AE",x"A5", -- 0x2648
    x"AF",x"49",x"FF",x"85",x"AF",x"A5",x"B9",x"49", -- 0x2650
    x"FF",x"85",x"B9",x"E6",x"B9",x"D0",x"0A",x"E6", -- 0x2658
    x"AF",x"D0",x"06",x"E6",x"AE",x"D0",x"02",x"E6", -- 0x2660
    x"AD",x"60",x"A2",x"0A",x"4C",x"2B",x"D1",x"A2", -- 0x2668
    x"74",x"B4",x"03",x"84",x"B9",x"B4",x"02",x"94", -- 0x2670
    x"03",x"B4",x"01",x"94",x"02",x"A4",x"B2",x"94", -- 0x2678
    x"01",x"69",x"08",x"30",x"EC",x"F0",x"EA",x"E9", -- 0x2680
    x"08",x"A8",x"A5",x"B9",x"B0",x"12",x"16",x"01", -- 0x2688
    x"90",x"02",x"F6",x"01",x"76",x"01",x"76",x"01", -- 0x2690
    x"76",x"02",x"76",x"03",x"6A",x"C8",x"D0",x"EE", -- 0x2698
    x"18",x"60",x"20",x"93",x"E8",x"F0",x"02",x"10", -- 0x26A0
    x"03",x"4C",x"D0",x"DE",x"A5",x"AC",x"E9",x"7F", -- 0x26A8
    x"48",x"A9",x"80",x"85",x"AC",x"A9",x"0F",x"A0", -- 0x26B0
    x"F1",x"20",x"65",x"E5",x"A9",x"13",x"A0",x"F1", -- 0x26B8
    x"20",x"A8",x"E7",x"A9",x"86",x"A0",x"F1",x"20", -- 0x26C0
    x"4A",x"E5",x"A9",x"02",x"A0",x"F1",x"20",x"FC", -- 0x26C8
    x"EB",x"A9",x"17",x"A0",x"F1",x"20",x"65",x"E5", -- 0x26D0
    x"68",x"20",x"F0",x"E9",x"A9",x"1B",x"A0",x"F1", -- 0x26D8
    x"20",x"32",x"E7",x"F0",x"4C",x"20",x"58",x"E7", -- 0x26E0
    x"A9",x"00",x"85",x"75",x"85",x"76",x"85",x"77", -- 0x26E8
    x"A5",x"B9",x"20",x"07",x"E7",x"A5",x"AF",x"20", -- 0x26F0
    x"07",x"E7",x"A5",x"AE",x"20",x"07",x"E7",x"A5", -- 0x26F8
    x"AD",x"20",x"0C",x"E7",x"4C",x"18",x"E8",x"D0", -- 0x2700
    x"03",x"4C",x"6F",x"E6",x"4A",x"09",x"80",x"A8", -- 0x2708
    x"90",x"13",x"18",x"A5",x"77",x"65",x"B6",x"85", -- 0x2710
    x"77",x"A5",x"76",x"65",x"B5",x"85",x"76",x"A5", -- 0x2718
    x"75",x"65",x"B4",x"85",x"75",x"66",x"75",x"66", -- 0x2720
    x"76",x"66",x"77",x"66",x"B9",x"98",x"4A",x"D0", -- 0x2728
    x"DE",x"60",x"85",x"71",x"84",x"72",x"A0",x"03", -- 0x2730
    x"B1",x"71",x"85",x"B6",x"88",x"B1",x"71",x"85", -- 0x2738
    x"B5",x"88",x"B1",x"71",x"85",x"B7",x"45",x"B0", -- 0x2740
    x"85",x"B8",x"A5",x"B7",x"09",x"80",x"85",x"B4", -- 0x2748
    x"88",x"B1",x"71",x"85",x"B3",x"A5",x"AC",x"60", -- 0x2750
    x"A5",x"B3",x"F0",x"1D",x"18",x"65",x"AC",x"90", -- 0x2758
    x"04",x"30",x"31",x"18",x"2C",x"10",x"12",x"69", -- 0x2760
    x"80",x"85",x"AC",x"D0",x"03",x"4C",x"FB",x"E5", -- 0x2768
    x"A5",x"B8",x"85",x"B0",x"60",x"A5",x"B0",x"10", -- 0x2770
    x"1B",x"68",x"68",x"4C",x"F7",x"E5",x"20",x"74", -- 0x2778
    x"E8",x"AA",x"F0",x"F0",x"18",x"69",x"02",x"B0", -- 0x2780
    x"0B",x"A2",x"00",x"86",x"B8",x"20",x"82",x"E5", -- 0x2788
    x"E6",x"AC",x"D0",x"E0",x"4C",x"6A",x"E6",x"20", -- 0x2790
    x"74",x"E8",x"A9",x"97",x"A0",x"F1",x"A2",x"00", -- 0x2798
    x"86",x"B8",x"20",x"27",x"E8",x"4C",x"AB",x"E7", -- 0x27A0
    x"20",x"32",x"E7",x"F0",x"66",x"20",x"83",x"E8", -- 0x27A8
    x"A9",x"00",x"38",x"E5",x"AC",x"85",x"AC",x"20", -- 0x27B0
    x"58",x"E7",x"E6",x"AC",x"F0",x"D6",x"A2",x"FD", -- 0x27B8
    x"A9",x"01",x"A4",x"B4",x"C4",x"AD",x"D0",x"0A", -- 0x27C0
    x"A4",x"B5",x"C4",x"AE",x"D0",x"04",x"A4",x"B6", -- 0x27C8
    x"C4",x"AF",x"08",x"2A",x"90",x"0A",x"E8",x"F0", -- 0x27D0
    x"2A",x"10",x"2C",x"A0",x"01",x"95",x"77",x"98", -- 0x27D8
    x"28",x"90",x"14",x"A8",x"A5",x"B6",x"E5",x"AF", -- 0x27E0
    x"85",x"B6",x"A5",x"B5",x"E5",x"AE",x"85",x"B5", -- 0x27E8
    x"A5",x"B4",x"E5",x"AD",x"85",x"B4",x"98",x"06", -- 0x27F0
    x"B6",x"26",x"B5",x"26",x"B4",x"B0",x"D3",x"30", -- 0x27F8
    x"C1",x"10",x"CF",x"A0",x"40",x"D0",x"D6",x"0A", -- 0x2800
    x"0A",x"0A",x"0A",x"0A",x"0A",x"85",x"B9",x"28", -- 0x2808
    x"4C",x"18",x"E8",x"A2",x"14",x"4C",x"2B",x"D1", -- 0x2810
    x"A5",x"75",x"85",x"AD",x"A5",x"76",x"85",x"AE", -- 0x2818
    x"A5",x"77",x"85",x"AF",x"4C",x"DB",x"E5",x"85", -- 0x2820
    x"71",x"84",x"72",x"A0",x"03",x"B1",x"71",x"85", -- 0x2828
    x"AF",x"88",x"B1",x"71",x"85",x"AE",x"88",x"B1", -- 0x2830
    x"71",x"85",x"B0",x"09",x"80",x"85",x"AD",x"88", -- 0x2838
    x"B1",x"71",x"85",x"AC",x"84",x"B9",x"60",x"A2", -- 0x2840
    x"A4",x"A0",x"00",x"F0",x"04",x"A6",x"97",x"A4", -- 0x2848
    x"98",x"20",x"83",x"E8",x"86",x"71",x"84",x"72", -- 0x2850
    x"A0",x"03",x"A5",x"AF",x"91",x"71",x"88",x"A5", -- 0x2858
    x"AE",x"91",x"71",x"88",x"A5",x"B0",x"09",x"7F", -- 0x2860
    x"25",x"AD",x"91",x"71",x"88",x"A5",x"AC",x"91", -- 0x2868
    x"71",x"84",x"B9",x"60",x"20",x"83",x"E8",x"A2", -- 0x2870
    x"05",x"B5",x"AB",x"95",x"B2",x"CA",x"D0",x"F9", -- 0x2878
    x"86",x"B9",x"60",x"A5",x"AC",x"F0",x"FB",x"06", -- 0x2880
    x"B9",x"90",x"F7",x"20",x"5F",x"E6",x"D0",x"F2", -- 0x2888
    x"4C",x"30",x"E6",x"A5",x"AC",x"F0",x"09",x"A5", -- 0x2890
    x"B0",x"2A",x"A9",x"FF",x"B0",x"02",x"A9",x"01", -- 0x2898
    x"60",x"20",x"93",x"E8",x"85",x"AD",x"A9",x"00", -- 0x28A0
    x"85",x"AE",x"A2",x"88",x"A5",x"AD",x"49",x"FF", -- 0x28A8
    x"2A",x"A9",x"00",x"85",x"AF",x"86",x"AC",x"85", -- 0x28B0
    x"B9",x"85",x"B0",x"4C",x"D6",x"E5",x"46",x"B0", -- 0x28B8
    x"60",x"85",x"73",x"84",x"74",x"A0",x"00",x"B1", -- 0x28C0
    x"73",x"C8",x"AA",x"F0",x"C6",x"B1",x"73",x"45", -- 0x28C8
    x"B0",x"30",x"C4",x"E4",x"AC",x"D0",x"1A",x"B1", -- 0x28D0
    x"73",x"09",x"80",x"C5",x"AD",x"D0",x"12",x"C8", -- 0x28D8
    x"B1",x"73",x"C5",x"AE",x"D0",x"0B",x"C8",x"A9", -- 0x28E0
    x"7F",x"C5",x"B9",x"B1",x"73",x"E5",x"AF",x"F0", -- 0x28E8
    x"28",x"A5",x"B0",x"90",x"02",x"49",x"FF",x"4C", -- 0x28F0
    x"99",x"E8",x"A5",x"AC",x"F0",x"4A",x"38",x"E9", -- 0x28F8
    x"98",x"24",x"B0",x"10",x"09",x"AA",x"A9",x"FF", -- 0x2900
    x"85",x"B2",x"20",x"43",x"E6",x"8A",x"A2",x"AC", -- 0x2908
    x"C9",x"F9",x"10",x"06",x"20",x"81",x"E6",x"84", -- 0x2910
    x"B2",x"60",x"A8",x"A5",x"B0",x"29",x"80",x"46", -- 0x2918
    x"AD",x"05",x"AD",x"85",x"AD",x"20",x"98",x"E6", -- 0x2920
    x"84",x"B2",x"60",x"A5",x"AC",x"C9",x"98",x"B0", -- 0x2928
    x"1E",x"20",x"FA",x"E8",x"84",x"B9",x"A5",x"B0", -- 0x2930
    x"84",x"B0",x"49",x"80",x"2A",x"A9",x"98",x"85", -- 0x2938
    x"AC",x"A5",x"AF",x"85",x"5B",x"4C",x"D6",x"E5", -- 0x2940
    x"85",x"AD",x"85",x"AE",x"85",x"AF",x"A8",x"60", -- 0x2948
    x"A0",x"00",x"84",x"5F",x"A2",x"09",x"94",x"A8", -- 0x2950
    x"CA",x"10",x"FB",x"90",x"7F",x"C9",x"2D",x"D0", -- 0x2958
    x"04",x"86",x"B1",x"F0",x"04",x"C9",x"2B",x"D0", -- 0x2960
    x"05",x"20",x"BC",x"00",x"90",x"6E",x"C9",x"24", -- 0x2968
    x"D0",x"03",x"4C",x"18",x"EE",x"C9",x"25",x"D0", -- 0x2970
    x"08",x"4C",x"46",x"EE",x"20",x"BC",x"00",x"90", -- 0x2978
    x"5B",x"C9",x"2E",x"F0",x"2E",x"C9",x"45",x"D0", -- 0x2980
    x"30",x"20",x"BC",x"00",x"90",x"17",x"C9",x"B6", -- 0x2988
    x"F0",x"0E",x"C9",x"2D",x"F0",x"0A",x"C9",x"B5", -- 0x2990
    x"F0",x"08",x"C9",x"2B",x"F0",x"04",x"D0",x"07", -- 0x2998
    x"66",x"AB",x"20",x"BC",x"00",x"90",x"5C",x"24", -- 0x29A0
    x"AB",x"10",x"0E",x"A9",x"00",x"38",x"E5",x"A9", -- 0x29A8
    x"4C",x"BB",x"E9",x"66",x"AA",x"24",x"AA",x"50", -- 0x29B0
    x"C3",x"A5",x"A9",x"38",x"E5",x"A8",x"85",x"A9", -- 0x29B8
    x"F0",x"12",x"10",x"09",x"20",x"97",x"E7",x"E6", -- 0x29C0
    x"A9",x"D0",x"F9",x"F0",x"07",x"20",x"7E",x"E7", -- 0x29C8
    x"C6",x"A9",x"D0",x"F9",x"A5",x"B1",x"30",x"01", -- 0x29D0
    x"60",x"4C",x"9F",x"EB",x"48",x"24",x"AA",x"10", -- 0x29D8
    x"02",x"E6",x"A8",x"20",x"7E",x"E7",x"68",x"38", -- 0x29E0
    x"E9",x"30",x"20",x"F0",x"E9",x"4C",x"7C",x"E9", -- 0x29E8
    x"48",x"20",x"74",x"E8",x"68",x"20",x"A4",x"E8", -- 0x29F0
    x"A5",x"B7",x"45",x"B0",x"85",x"B8",x"A6",x"AC", -- 0x29F8
    x"4C",x"68",x"E5",x"A5",x"A9",x"C9",x"0A",x"90", -- 0x2A00
    x"09",x"A9",x"64",x"24",x"AB",x"30",x"0E",x"4C", -- 0x2A08
    x"6A",x"E6",x"0A",x"0A",x"65",x"A9",x"0A",x"A0", -- 0x2A10
    x"00",x"71",x"C3",x"E9",x"2F",x"85",x"A9",x"4C", -- 0x2A18
    x"A2",x"E9",x"A9",x"8B",x"A0",x"F7",x"20",x"7A", -- 0x2A20
    x"D8",x"A5",x"88",x"A6",x"87",x"85",x"AD",x"86", -- 0x2A28
    x"AE",x"A2",x"90",x"38",x"20",x"B1",x"E8",x"A0", -- 0x2A30
    x"00",x"98",x"20",x"4D",x"EA",x"4C",x"7A",x"D8", -- 0x2A38
    x"A0",x"01",x"A9",x"20",x"24",x"B0",x"10",x"02", -- 0x2A40
    x"A9",x"2D",x"99",x"EF",x"00",x"85",x"B0",x"84", -- 0x2A48
    x"BA",x"C8",x"A6",x"AC",x"D0",x"05",x"A9",x"30", -- 0x2A50
    x"4C",x"59",x"EB",x"A9",x"00",x"E0",x"81",x"B0", -- 0x2A58
    x"09",x"A9",x"27",x"A0",x"F1",x"20",x"E0",x"E6", -- 0x2A60
    x"A9",x"FA",x"85",x"A8",x"A9",x"23",x"A0",x"F1", -- 0x2A68
    x"20",x"C1",x"E8",x"F0",x"1E",x"10",x"12",x"A9", -- 0x2A70
    x"1F",x"A0",x"F1",x"20",x"C1",x"E8",x"F0",x"02", -- 0x2A78
    x"10",x"0E",x"20",x"7E",x"E7",x"C6",x"A8",x"D0", -- 0x2A80
    x"EE",x"20",x"97",x"E7",x"E6",x"A8",x"D0",x"DC", -- 0x2A88
    x"20",x"61",x"E5",x"20",x"FA",x"E8",x"A2",x"01", -- 0x2A90
    x"A5",x"A8",x"18",x"69",x"07",x"30",x"09",x"C9", -- 0x2A98
    x"08",x"B0",x"06",x"69",x"FF",x"AA",x"A9",x"02", -- 0x2AA0
    x"38",x"E9",x"02",x"85",x"A9",x"86",x"A8",x"8A", -- 0x2AA8
    x"F0",x"02",x"10",x"13",x"A4",x"BA",x"A9",x"2E", -- 0x2AB0
    x"C8",x"99",x"EF",x"00",x"8A",x"F0",x"06",x"A9", -- 0x2AB8
    x"30",x"C8",x"99",x"EF",x"00",x"84",x"BA",x"A0", -- 0x2AC0
    x"00",x"A2",x"80",x"A5",x"AF",x"18",x"79",x"9D", -- 0x2AC8
    x"F1",x"85",x"AF",x"A5",x"AE",x"79",x"9C",x"F1", -- 0x2AD0
    x"85",x"AE",x"A5",x"AD",x"79",x"9B",x"F1",x"85", -- 0x2AD8
    x"AD",x"E8",x"B0",x"04",x"10",x"E5",x"30",x"02", -- 0x2AE0
    x"30",x"E1",x"8A",x"90",x"04",x"49",x"FF",x"69", -- 0x2AE8
    x"0A",x"69",x"2F",x"C8",x"C8",x"C8",x"84",x"95", -- 0x2AF0
    x"A4",x"BA",x"C8",x"AA",x"29",x"7F",x"99",x"EF", -- 0x2AF8
    x"00",x"C6",x"A8",x"D0",x"06",x"A9",x"2E",x"C8", -- 0x2B00
    x"99",x"EF",x"00",x"84",x"BA",x"A4",x"95",x"8A", -- 0x2B08
    x"49",x"FF",x"29",x"80",x"AA",x"C0",x"12",x"D0", -- 0x2B10
    x"B2",x"A4",x"BA",x"B9",x"EF",x"00",x"88",x"C9", -- 0x2B18
    x"30",x"F0",x"F8",x"C9",x"2E",x"F0",x"01",x"C8", -- 0x2B20
    x"A9",x"2B",x"A6",x"A9",x"F0",x"2E",x"10",x"08", -- 0x2B28
    x"A9",x"00",x"38",x"E5",x"A9",x"AA",x"A9",x"2D", -- 0x2B30
    x"99",x"F1",x"00",x"A9",x"45",x"99",x"F0",x"00", -- 0x2B38
    x"8A",x"A2",x"2F",x"38",x"E8",x"E9",x"0A",x"B0", -- 0x2B40
    x"FB",x"69",x"3A",x"99",x"F3",x"00",x"8A",x"99", -- 0x2B48
    x"F2",x"00",x"A9",x"00",x"99",x"F4",x"00",x"F0", -- 0x2B50
    x"08",x"99",x"EF",x"00",x"A9",x"00",x"99",x"F0", -- 0x2B58
    x"00",x"A9",x"F0",x"A0",x"00",x"60",x"F0",x"42", -- 0x2B60
    x"A5",x"B3",x"D0",x"03",x"4C",x"F9",x"E5",x"A2", -- 0x2B68
    x"9C",x"A0",x"00",x"20",x"51",x"E8",x"A5",x"B7", -- 0x2B70
    x"10",x"0F",x"20",x"2B",x"E9",x"A9",x"9C",x"A0", -- 0x2B78
    x"00",x"20",x"C1",x"E8",x"D0",x"03",x"98",x"A4", -- 0x2B80
    x"5B",x"20",x"6C",x"E5",x"98",x"48",x"20",x"A2", -- 0x2B88
    x"E6",x"A9",x"9C",x"A0",x"00",x"20",x"E0",x"E6", -- 0x2B90
    x"20",x"AA",x"EB",x"68",x"4A",x"90",x"0A",x"A5", -- 0x2B98
    x"AC",x"F0",x"06",x"A5",x"B0",x"49",x"FF",x"85", -- 0x2BA0
    x"B0",x"60",x"A9",x"2B",x"A0",x"F1",x"20",x"E0", -- 0x2BA8
    x"E6",x"A5",x"B9",x"69",x"50",x"90",x"03",x"20", -- 0x2BB0
    x"8B",x"E8",x"85",x"A3",x"20",x"77",x"E8",x"A5", -- 0x2BB8
    x"AC",x"C9",x"88",x"90",x"03",x"20",x"75",x"E7", -- 0x2BC0
    x"20",x"2B",x"E9",x"A5",x"5B",x"18",x"69",x"81", -- 0x2BC8
    x"F0",x"F3",x"38",x"E9",x"01",x"48",x"A2",x"04", -- 0x2BD0
    x"B5",x"B3",x"B4",x"AC",x"95",x"AC",x"94",x"B3", -- 0x2BD8
    x"CA",x"10",x"F5",x"A5",x"A3",x"85",x"B9",x"20", -- 0x2BE0
    x"4D",x"E5",x"20",x"9F",x"EB",x"A9",x"2F",x"A0", -- 0x2BE8
    x"F1",x"20",x"12",x"EC",x"A9",x"00",x"85",x"B8", -- 0x2BF0
    x"68",x"4C",x"5A",x"E7",x"85",x"BA",x"84",x"BB", -- 0x2BF8
    x"20",x"47",x"E8",x"A9",x"A4",x"20",x"E0",x"E6", -- 0x2C00
    x"20",x"16",x"EC",x"A9",x"A4",x"A0",x"00",x"4C", -- 0x2C08
    x"E0",x"E6",x"85",x"BA",x"84",x"BB",x"A2",x"A8", -- 0x2C10
    x"20",x"49",x"E8",x"B1",x"BA",x"85",x"B1",x"A4", -- 0x2C18
    x"BA",x"C8",x"98",x"D0",x"02",x"E6",x"BB",x"85", -- 0x2C20
    x"BA",x"A4",x"BB",x"20",x"E0",x"E6",x"A5",x"BA", -- 0x2C28
    x"A4",x"BB",x"18",x"69",x"04",x"90",x"01",x"C8", -- 0x2C30
    x"85",x"BA",x"84",x"BB",x"20",x"65",x"E5",x"A9", -- 0x2C38
    x"A8",x"A0",x"00",x"C6",x"B1",x"D0",x"E4",x"60", -- 0x2C40
    x"A5",x"AC",x"F0",x"07",x"A2",x"D4",x"A0",x"00", -- 0x2C48
    x"20",x"51",x"E8",x"A0",x"13",x"06",x"D7",x"26", -- 0x2C50
    x"D6",x"26",x"D5",x"26",x"D4",x"90",x"06",x"A9", -- 0x2C58
    x"AF",x"45",x"D7",x"85",x"D7",x"88",x"D0",x"ED", -- 0x2C60
    x"A2",x"02",x"B5",x"D4",x"95",x"AD",x"CA",x"10", -- 0x2C68
    x"F9",x"A9",x"80",x"85",x"AC",x"0A",x"85",x"B0", -- 0x2C70
    x"4C",x"DB",x"E5",x"A9",x"4C",x"A0",x"F1",x"20", -- 0x2C78
    x"65",x"E5",x"20",x"74",x"E8",x"A9",x"61",x"A0", -- 0x2C80
    x"F1",x"A6",x"B7",x"20",x"A0",x"E7",x"20",x"74", -- 0x2C88
    x"E8",x"20",x"2B",x"E9",x"A9",x"00",x"85",x"B8", -- 0x2C90
    x"20",x"4D",x"E5",x"A9",x"93",x"A0",x"F1",x"20", -- 0x2C98
    x"4A",x"E5",x"A5",x"B0",x"48",x"10",x"0D",x"20", -- 0x2CA0
    x"61",x"E5",x"A5",x"B0",x"30",x"09",x"A5",x"63", -- 0x2CA8
    x"49",x"FF",x"85",x"63",x"20",x"9F",x"EB",x"A9", -- 0x2CB0
    x"93",x"A0",x"F1",x"20",x"65",x"E5",x"68",x"10", -- 0x2CB8
    x"03",x"20",x"9F",x"EB",x"A9",x"50",x"A0",x"F1", -- 0x2CC0
    x"4C",x"FC",x"EB",x"20",x"47",x"E8",x"A9",x"00", -- 0x2CC8
    x"85",x"63",x"20",x"82",x"EC",x"A2",x"9C",x"A0", -- 0x2CD0
    x"00",x"20",x"51",x"E8",x"A9",x"A4",x"A0",x"00", -- 0x2CD8
    x"20",x"27",x"E8",x"A9",x"00",x"85",x"B0",x"A5", -- 0x2CE0
    x"63",x"20",x"F3",x"EC",x"A9",x"9C",x"A0",x"00", -- 0x2CE8
    x"4C",x"A8",x"E7",x"48",x"4C",x"B4",x"EC",x"20", -- 0x2CF0
    x"0A",x"00",x"4C",x"96",x"DB",x"A5",x"B0",x"48", -- 0x2CF8
    x"10",x"03",x"20",x"9F",x"EB",x"A5",x"AC",x"48", -- 0x2D00
    x"C9",x"81",x"90",x"07",x"A9",x"86",x"A0",x"F1", -- 0x2D08
    x"20",x"A8",x"E7",x"A9",x"65",x"A0",x"F1",x"20", -- 0x2D10
    x"FC",x"EB",x"68",x"C9",x"81",x"90",x"07",x"A9", -- 0x2D18
    x"4C",x"A0",x"F1",x"20",x"4A",x"E5",x"68",x"10", -- 0x2D20
    x"16",x"4C",x"9F",x"EB",x"20",x"7F",x"E4",x"E0", -- 0x2D28
    x"08",x"B0",x"20",x"A9",x"00",x"38",x"2A",x"CA", -- 0x2D30
    x"10",x"FC",x"E8",x"01",x"11",x"81",x"11",x"60", -- 0x2D38
    x"20",x"7F",x"E4",x"E0",x"08",x"B0",x"0C",x"A9", -- 0x2D40
    x"FF",x"2A",x"CA",x"10",x"FC",x"E8",x"21",x"11", -- 0x2D48
    x"81",x"11",x"60",x"4C",x"D0",x"DE",x"20",x"BC", -- 0x2D50
    x"00",x"20",x"7F",x"E4",x"E0",x"08",x"B0",x"F3", -- 0x2D58
    x"20",x"C2",x"00",x"C9",x"29",x"F0",x"03",x"4C", -- 0x2D60
    x"A9",x"DB",x"20",x"BC",x"00",x"A9",x"00",x"38", -- 0x2D68
    x"2A",x"CA",x"10",x"FC",x"E8",x"21",x"11",x"F0", -- 0x2D70
    x"02",x"A9",x"FF",x"4C",x"A4",x"E8",x"E0",x"19", -- 0x2D78
    x"B0",x"48",x"86",x"78",x"A9",x"18",x"20",x"E1", -- 0x2D80
    x"E0",x"A0",x"17",x"A2",x"18",x"46",x"11",x"66", -- 0x2D88
    x"12",x"66",x"13",x"8A",x"2A",x"91",x"AD",x"88", -- 0x2D90
    x"10",x"F3",x"A5",x"78",x"F0",x"0A",x"AA",x"38", -- 0x2D98
    x"49",x"FF",x"69",x"18",x"F0",x"1C",x"D0",x"0F", -- 0x2DA0
    x"A8",x"B1",x"AD",x"C9",x"30",x"D0",x"07",x"CA", -- 0x2DA8
    x"F0",x"03",x"C8",x"10",x"F4",x"E8",x"98",x"18", -- 0x2DB0
    x"65",x"AD",x"85",x"AD",x"A9",x"00",x"65",x"AE", -- 0x2DB8
    x"85",x"AE",x"86",x"AC",x"20",x"BC",x"00",x"4C", -- 0x2DC0
    x"2C",x"E1",x"4C",x"D0",x"DE",x"E0",x"07",x"B0", -- 0x2DC8
    x"F9",x"86",x"78",x"A9",x"06",x"20",x"E1",x"E0", -- 0x2DD0
    x"A0",x"05",x"F8",x"A5",x"13",x"20",x"FB",x"ED", -- 0x2DD8
    x"A5",x"12",x"20",x"FB",x"ED",x"A5",x"11",x"20", -- 0x2DE0
    x"FB",x"ED",x"D8",x"A2",x"06",x"A5",x"78",x"F0", -- 0x2DE8
    x"B7",x"AA",x"38",x"49",x"FF",x"69",x"06",x"F0", -- 0x2DF0
    x"C9",x"D0",x"BC",x"AA",x"29",x"0F",x"20",x"06", -- 0x2DF8
    x"EE",x"8A",x"4A",x"4A",x"4A",x"4A",x"C9",x"0A", -- 0x2E00
    x"69",x"30",x"91",x"AD",x"88",x"60",x"85",x"AC", -- 0x2E08
    x"A9",x"00",x"85",x"B8",x"8A",x"20",x"F0",x"E9", -- 0x2E10
    x"20",x"BC",x"00",x"90",x"0A",x"09",x"20",x"E9", -- 0x2E18
    x"61",x"C9",x"06",x"B0",x"2A",x"69",x"0A",x"29", -- 0x2E20
    x"0F",x"AA",x"A5",x"AC",x"F0",x"E4",x"69",x"04", -- 0x2E28
    x"90",x"DC",x"4C",x"6A",x"E6",x"AA",x"A5",x"AC", -- 0x2E30
    x"F0",x"06",x"E6",x"AC",x"F0",x"F4",x"A9",x"00", -- 0x2E38
    x"85",x"B8",x"8A",x"20",x"F0",x"E9",x"20",x"BC", -- 0x2E40
    x"00",x"49",x"30",x"C9",x"02",x"90",x"E6",x"4C", -- 0x2E48
    x"D4",x"E9",x"AD",x"00",x"02",x"D0",x"18",x"20", -- 0x2E50
    x"94",x"F0",x"90",x"0B",x"8D",x"01",x"02",x"A2", -- 0x2E58
    x"20",x"8E",x"02",x"02",x"4C",x"06",x"D5",x"AE", -- 0x2E60
    x"02",x"02",x"F0",x"03",x"CE",x"02",x"02",x"A2", -- 0x2E68
    x"D8",x"20",x"7A",x"EE",x"A2",x"DB",x"20",x"7A", -- 0x2E70
    x"EE",x"60",x"B5",x"00",x"10",x"FB",x"0A",x"29", -- 0x2E78
    x"40",x"F0",x"F6",x"95",x"00",x"8A",x"A8",x"68", -- 0x2E80
    x"68",x"A9",x"05",x"20",x"F4",x"D0",x"A5",x"C4", -- 0x2E88
    x"48",x"A5",x"C3",x"48",x"A5",x"88",x"48",x"A5", -- 0x2E90
    x"87",x"48",x"A9",x"8D",x"48",x"B9",x"01",x"00", -- 0x2E98
    x"85",x"C3",x"B9",x"02",x"00",x"85",x"C4",x"4C", -- 0x2EA0
    x"AB",x"D4",x"20",x"94",x"F0",x"B0",x"09",x"AD", -- 0x2EA8
    x"02",x"02",x"F0",x"09",x"AD",x"01",x"02",x"38", -- 0x2EB0
    x"A2",x"00",x"8E",x"02",x"02",x"60",x"A2",x"DB", -- 0x2EB8
    x"2C",x"A2",x"D8",x"C9",x"93",x"F0",x"11",x"C9", -- 0x2EC0
    x"B4",x"F0",x"07",x"49",x"A2",x"F0",x"0E",x"4C", -- 0x2EC8
    x"A9",x"DB",x"A9",x"7F",x"35",x"00",x"10",x"05", -- 0x2ED0
    x"B5",x"00",x"0A",x"15",x"00",x"95",x"00",x"4C", -- 0x2ED8
    x"BC",x"00",x"58",x"A2",x"DB",x"2C",x"A2",x"D8", -- 0x2EE0
    x"86",x"78",x"20",x"BC",x"00",x"20",x"FA",x"D6", -- 0x2EE8
    x"A5",x"79",x"A6",x"7A",x"20",x"17",x"D3",x"B0", -- 0x2EF0
    x"03",x"4C",x"61",x"D6",x"A6",x"78",x"A5",x"AA", -- 0x2EF8
    x"E9",x"01",x"95",x"01",x"A5",x"AB",x"E9",x"00", -- 0x2F00
    x"95",x"02",x"A9",x"C0",x"95",x"00",x"60",x"D0", -- 0x2F08
    x"FD",x"A5",x"DB",x"0A",x"05",x"DB",x"85",x"DB", -- 0x2F10
    x"4C",x"68",x"D6",x"D0",x"F1",x"A5",x"D8",x"0A", -- 0x2F18
    x"05",x"D8",x"85",x"D8",x"4C",x"68",x"D6",x"20", -- 0x2F20
    x"90",x"DA",x"4C",x"77",x"DA",x"20",x"5B",x"EF", -- 0x2F28
    x"10",x"FB",x"A5",x"B4",x"09",x"80",x"85",x"B4", -- 0x2F30
    x"20",x"6A",x"E5",x"F0",x"F0",x"20",x"5B",x"EF", -- 0x2F38
    x"30",x"FB",x"F0",x"F9",x"A5",x"B4",x"09",x"80", -- 0x2F40
    x"85",x"B4",x"20",x"6A",x"E5",x"F0",x"EE",x"C9", -- 0x2F48
    x"29",x"D0",x"05",x"68",x"68",x"4C",x"BC",x"00", -- 0x2F50
    x"4C",x"A9",x"DB",x"20",x"C2",x"00",x"C9",x"2C", -- 0x2F58
    x"D0",x"ED",x"20",x"83",x"E8",x"A5",x"B0",x"09", -- 0x2F60
    x"7F",x"25",x"AD",x"48",x"A5",x"AE",x"48",x"A5", -- 0x2F68
    x"AF",x"48",x"A5",x"AC",x"48",x"20",x"BC",x"00", -- 0x2F70
    x"20",x"74",x"DA",x"68",x"85",x"B3",x"68",x"85", -- 0x2F78
    x"B6",x"68",x"85",x"B5",x"68",x"85",x"B4",x"85", -- 0x2F80
    x"B7",x"A9",x"B3",x"A0",x"00",x"4C",x"C1",x"E8", -- 0x2F88
    x"C9",x"2C",x"F0",x"1B",x"20",x"33",x"E4",x"8A", -- 0x2F90
    x"F0",x"0A",x"E0",x"10",x"90",x"45",x"E4",x"64", -- 0x2F98
    x"B0",x"02",x"86",x"64",x"86",x"0F",x"20",x"C2", -- 0x2FA0
    x"00",x"F0",x"1A",x"C9",x"2C",x"D0",x"A9",x"20", -- 0x2FA8
    x"30",x"E4",x"8A",x"30",x"2E",x"E0",x"01",x"90", -- 0x2FB0
    x"2A",x"A5",x"0F",x"F0",x"06",x"E4",x"0F",x"F0", -- 0x2FB8
    x"02",x"B0",x"20",x"86",x"64",x"A5",x"0F",x"F0", -- 0x2FC0
    x"06",x"C5",x"64",x"B0",x"03",x"85",x"64",x"38", -- 0x2FC8
    x"E5",x"64",x"B0",x"FC",x"65",x"64",x"18",x"65", -- 0x2FD0
    x"64",x"85",x"10",x"A5",x"0F",x"38",x"E5",x"10", -- 0x2FD8
    x"85",x"10",x"60",x"4C",x"D0",x"DE",x"A5",x"B0", -- 0x2FE0
    x"30",x"F9",x"A5",x"AC",x"F0",x"F4",x"20",x"74", -- 0x2FE8
    x"E8",x"A9",x"00",x"85",x"77",x"85",x"76",x"85", -- 0x2FF0
    x"75",x"85",x"78",x"85",x"AF",x"85",x"AE",x"85", -- 0x2FF8
    x"AD",x"A2",x"18",x"A5",x"B3",x"4A",x"B0",x"0E", -- 0x3000
    x"06",x"B6",x"26",x"B5",x"26",x"B4",x"26",x"77", -- 0x3008
    x"26",x"76",x"26",x"75",x"26",x"78",x"06",x"B6", -- 0x3010
    x"26",x"B5",x"26",x"B4",x"26",x"77",x"26",x"76", -- 0x3018
    x"26",x"75",x"26",x"78",x"06",x"AF",x"26",x"AE", -- 0x3020
    x"26",x"AD",x"A5",x"AF",x"2A",x"85",x"5B",x"A5", -- 0x3028
    x"AE",x"2A",x"85",x"5C",x"A5",x"AD",x"2A",x"85", -- 0x3030
    x"5D",x"A9",x"00",x"2A",x"85",x"5E",x"A5",x"77", -- 0x3038
    x"E5",x"5B",x"85",x"5B",x"A5",x"76",x"E5",x"5C", -- 0x3040
    x"85",x"5C",x"A5",x"75",x"E5",x"5D",x"A8",x"A5", -- 0x3048
    x"78",x"E5",x"5E",x"90",x"0E",x"85",x"78",x"84", -- 0x3050
    x"75",x"A5",x"5C",x"85",x"76",x"A5",x"5B",x"85", -- 0x3058
    x"77",x"E6",x"AF",x"CA",x"D0",x"A2",x"38",x"A5", -- 0x3060
    x"B3",x"E9",x"80",x"6A",x"69",x"00",x"85",x"AC", -- 0x3068
    x"4C",x"DB",x"E5",x"20",x"BC",x"00",x"20",x"51", -- 0x3070
    x"DD",x"20",x"96",x"DB",x"A4",x"95",x"A5",x"96", -- 0x3078
    x"4C",x"00",x"E0",x"A9",x"61",x"A0",x"F1",x"20", -- 0x3080
    x"27",x"E8",x"C6",x"AC",x"60",x"A9",x"61",x"A0", -- 0x3088
    x"F1",x"4C",x"27",x"E8",x"6C",x"05",x"02",x"6C", -- 0x3090
    x"07",x"02",x"6C",x"09",x"02",x"6C",x"0B",x"02", -- 0x3098
    x"00",x"00",x"00",x"52",x"EE",x"E6",x"C3",x"D0", -- 0x30A0
    x"02",x"E6",x"C4",x"AD",x"FF",x"FF",x"C9",x"3A", -- 0x30A8
    x"B0",x"0A",x"C9",x"20",x"F0",x"EF",x"38",x"E9", -- 0x30B0
    x"30",x"38",x"E9",x"D0",x"60",x"4C",x"00",x"D0", -- 0x30B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4C", -- 0x30C0
    x"D0",x"DE",x"00",x"00",x"00",x"F2",x"00",x"04", -- 0x30C8
    x"0D",x"0A",x"4D",x"65",x"6D",x"6F",x"72",x"79", -- 0x30D0
    x"20",x"73",x"69",x"7A",x"65",x"20",x"00",x"20", -- 0x30D8
    x"42",x"79",x"74",x"65",x"73",x"20",x"66",x"72", -- 0x30E0
    x"65",x"65",x"0D",x"0A",x"0A",x"45",x"6E",x"68", -- 0x30E8
    x"61",x"6E",x"63",x"65",x"64",x"20",x"42",x"41", -- 0x30F0
    x"53",x"49",x"43",x"20",x"32",x"2E",x"30",x"39", -- 0x30F8
    x"0A",x"00",x"02",x"80",x"19",x"56",x"62",x"80", -- 0x3100
    x"76",x"22",x"F3",x"82",x"38",x"AA",x"40",x"80", -- 0x3108
    x"35",x"04",x"F3",x"81",x"35",x"04",x"F3",x"80", -- 0x3110
    x"80",x"00",x"00",x"80",x"31",x"72",x"18",x"91", -- 0x3118
    x"43",x"4F",x"F8",x"94",x"74",x"23",x"F7",x"94", -- 0x3120
    x"74",x"24",x"00",x"81",x"38",x"AA",x"3B",x"06", -- 0x3128
    x"74",x"63",x"90",x"8C",x"77",x"23",x"0C",x"AB", -- 0x3130
    x"7A",x"1E",x"94",x"00",x"7C",x"63",x"42",x"80", -- 0x3138
    x"7E",x"75",x"FE",x"D0",x"80",x"31",x"72",x"15", -- 0x3140
    x"81",x"00",x"00",x"00",x"81",x"49",x"0F",x"DB", -- 0x3148
    x"04",x"86",x"1E",x"D7",x"FB",x"87",x"99",x"26", -- 0x3150
    x"65",x"87",x"23",x"34",x"58",x"86",x"A5",x"5D", -- 0x3158
    x"E1",x"83",x"49",x"0F",x"DB",x"08",x"78",x"3A", -- 0x3160
    x"C5",x"37",x"7B",x"83",x"A2",x"5C",x"7C",x"2E", -- 0x3168
    x"DD",x"4D",x"7D",x"99",x"B0",x"1E",x"7D",x"59", -- 0x3170
    x"ED",x"24",x"7E",x"91",x"72",x"00",x"7E",x"4C", -- 0x3178
    x"B9",x"73",x"7F",x"AA",x"AA",x"53",x"81",x"00", -- 0x3180
    x"00",x"00",x"81",x"80",x"00",x"00",x"90",x"80", -- 0x3188
    x"00",x"00",x"00",x"7F",x"00",x"00",x"00",x"84", -- 0x3190
    x"20",x"00",x"00",x"FE",x"79",x"60",x"00",x"27", -- 0x3198
    x"10",x"FF",x"FC",x"18",x"00",x"00",x"64",x"FF", -- 0x31A0
    x"FF",x"F6",x"00",x"00",x"01",x"09",x"D5",x"46", -- 0x31A8
    x"D4",x"0B",x"DA",x"7A",x"D6",x"ED",x"D8",x"05", -- 0x31B0
    x"DD",x"0D",x"D9",x"58",x"D7",x"2A",x"D7",x"D9", -- 0x31B8
    x"D5",x"98",x"D5",x"A8",x"D6",x"30",x"D5",x"BC", -- 0x31C0
    x"D5",x"0E",x"EF",x"1A",x"EF",x"65",x"D6",x"BB", -- 0x31C8
    x"D6",x"07",x"D5",x"CB",x"D6",x"6E",x"D5",x"2D", -- 0x31D0
    x"D7",x"2F",x"E5",x"99",x"F0",x"9C",x"F0",x"1A", -- 0x31D8
    x"E0",x"B4",x"E4",x"D0",x"E4",x"1D",x"E5",x"A2", -- 0x31E0
    x"D5",x"0B",x"D6",x"F9",x"D7",x"74",x"D5",x"91", -- 0x31E8
    x"D3",x"8E",x"D3",x"3C",x"D3",x"8F",x"EF",x"C8", -- 0x31F0
    x"D7",x"F5",x"E4",x"2B",x"ED",x"3F",x"ED",x"BD", -- 0x31F8
    x"EE",x"C0",x"EE",x"0B",x"DC",x"0B",x"DC",x"0B", -- 0x3200
    x"DC",x"8F",x"DA",x"92",x"DB",x"92",x"DB",x"0B", -- 0x3208
    x"DC",x"0B",x"DC",x"0B",x"DC",x"0B",x"DC",x"0B", -- 0x3210
    x"DC",x"0B",x"DC",x"0B",x"DC",x"0B",x"DC",x"0B", -- 0x3218
    x"DC",x"0B",x"DC",x"00",x"00",x"05",x"DC",x"0B", -- 0x3220
    x"DC",x"05",x"DC",x"05",x"DC",x"05",x"DC",x"05", -- 0x3228
    x"DC",x"0B",x"DC",x"32",x"DC",x"32",x"DC",x"00", -- 0x3230
    x"00",x"26",x"EF",x"26",x"EF",x"11",x"DC",x"11", -- 0x3238
    x"DC",x"00",x"00",x"16",x"DC",x"16",x"DC",x"16", -- 0x3240
    x"DC",x"A0",x"E8",x"2A",x"E9",x"BD",x"E8",x"F6", -- 0x3248
    x"EC",x"EB",x"DF",x"0A",x"E0",x"E5",x"EF",x"47", -- 0x3250
    x"EC",x"A1",x"E6",x"A9",x"EB",x"7A",x"EC",x"81", -- 0x3258
    x"EC",x"CA",x"EC",x"FC",x"EC",x"A9",x"E4",x"BD", -- 0x3260
    x"E4",x"FB",x"E3",x"14",x"E4",x"CC",x"E0",x"41", -- 0x3268
    x"E4",x"1F",x"E4",x"D9",x"E3",x"B8",x"E3",x"2A", -- 0x3270
    x"E3",x"CC",x"ED",x"7D",x"ED",x"55",x"ED",x"2C", -- 0x3278
    x"EF",x"3C",x"EF",x"82",x"F0",x"8C",x"F0",x"72", -- 0x3280
    x"F0",x"3C",x"E3",x"45",x"E3",x"74",x"E3",x"79", -- 0x3288
    x"67",x"E5",x"79",x"4C",x"E5",x"7B",x"E2",x"E6", -- 0x3290
    x"7B",x"AA",x"E7",x"7F",x"65",x"EB",x"50",x"7B", -- 0x3298
    x"DC",x"46",x"61",x"DC",x"46",x"6E",x"DC",x"56", -- 0x32A0
    x"27",x"DD",x"56",x"0F",x"DD",x"7D",x"9E",x"EB", -- 0x32A8
    x"5A",x"BD",x"DB",x"64",x"9C",x"DC",x"2A",x"2B", -- 0x32B0
    x"2D",x"2F",x"3C",x"3D",x"3E",x"3F",x"41",x"42", -- 0x32B8
    x"43",x"44",x"45",x"46",x"47",x"48",x"49",x"4C", -- 0x32C0
    x"4D",x"4E",x"4F",x"50",x"52",x"53",x"54",x"55", -- 0x32C8
    x"56",x"57",x"5E",x"00",x"0E",x"F3",x"10",x"F3", -- 0x32D0
    x"12",x"F3",x"14",x"F3",x"16",x"F3",x"1A",x"F3", -- 0x32D8
    x"1C",x"F3",x"20",x"F3",x"22",x"F3",x"32",x"F3", -- 0x32E0
    x"4B",x"F3",x"62",x"F3",x"7B",x"F3",x"86",x"F3", -- 0x32E8
    x"90",x"F3",x"9D",x"F3",x"A3",x"F3",x"B5",x"F3", -- 0x32F0
    x"DA",x"F3",x"E8",x"F3",x"FA",x"F3",x"02",x"F4", -- 0x32F8
    x"17",x"F4",x"46",x"F4",x"71",x"F4",x"85",x"F4", -- 0x3300
    x"96",x"F4",x"A2",x"F4",x"B1",x"F4",x"B7",x"00", -- 0x3308
    x"B5",x"00",x"B6",x"00",x"B8",x"00",x"3C",x"BE", -- 0x3310
    x"C1",x"00",x"C0",x"00",x"3E",x"BD",x"BF",x"00", -- 0x3318
    x"9F",x"00",x"42",x"53",x"28",x"C4",x"4E",x"44", -- 0x3320
    x"BA",x"53",x"43",x"28",x"D6",x"54",x"4E",x"28", -- 0x3328
    x"CF",x"00",x"49",x"4E",x"24",x"28",x"DB",x"49", -- 0x3330
    x"54",x"43",x"4C",x"52",x"A8",x"49",x"54",x"53", -- 0x3338
    x"45",x"54",x"A7",x"49",x"54",x"54",x"53",x"54", -- 0x3340
    x"28",x"DC",x"00",x"41",x"4C",x"4C",x"9C",x"48", -- 0x3348
    x"52",x"24",x"28",x"D9",x"4C",x"45",x"41",x"52", -- 0x3350
    x"A2",x"4F",x"4E",x"54",x"A0",x"4F",x"53",x"28", -- 0x3358
    x"CC",x"00",x"41",x"54",x"41",x"83",x"45",x"43", -- 0x3360
    x"88",x"45",x"45",x"4B",x"28",x"D1",x"45",x"46", -- 0x3368
    x"99",x"49",x"4D",x"85",x"4F",x"4B",x"45",x"9B", -- 0x3370
    x"4F",x"9D",x"00",x"4E",x"44",x"80",x"4F",x"52", -- 0x3378
    x"BB",x"58",x"50",x"28",x"CB",x"00",x"4E",x"AD", -- 0x3380
    x"4F",x"52",x"81",x"52",x"45",x"28",x"C6",x"00", -- 0x3388
    x"45",x"54",x"A5",x"4F",x"53",x"55",x"42",x"8D", -- 0x3390
    x"4F",x"54",x"4F",x"89",x"00",x"45",x"58",x"24", -- 0x3398
    x"28",x"DA",x"00",x"46",x"8B",x"4E",x"43",x"95", -- 0x33A0
    x"4E",x"50",x"55",x"54",x"84",x"4E",x"54",x"28", -- 0x33A8
    x"C3",x"52",x"51",x"A9",x"00",x"43",x"41",x"53", -- 0x33B0
    x"45",x"24",x"28",x"D8",x"45",x"46",x"54",x"24", -- 0x33B8
    x"28",x"E2",x"45",x"4E",x"28",x"D3",x"45",x"54", -- 0x33C0
    x"87",x"49",x"53",x"54",x"A1",x"4F",x"41",x"44", -- 0x33C8
    x"97",x"4F",x"47",x"28",x"CA",x"4F",x"4F",x"50", -- 0x33D0
    x"9E",x"00",x"41",x"58",x"28",x"DD",x"49",x"44", -- 0x33D8
    x"24",x"28",x"E4",x"49",x"4E",x"28",x"DE",x"00", -- 0x33E0
    x"45",x"57",x"A3",x"45",x"58",x"54",x"82",x"4D", -- 0x33E8
    x"49",x"AA",x"4F",x"54",x"B0",x"55",x"4C",x"4C", -- 0x33F0
    x"94",x"00",x"46",x"46",x"B4",x"4E",x"93",x"52", -- 0x33F8
    x"BC",x"00",x"45",x"45",x"4B",x"28",x"D0",x"49", -- 0x3400
    x"DF",x"4F",x"4B",x"45",x"9A",x"4F",x"53",x"28", -- 0x3408
    x"C7",x"52",x"49",x"4E",x"54",x"9F",x"00",x"45", -- 0x3410
    x"41",x"44",x"86",x"45",x"4D",x"91",x"45",x"53", -- 0x3418
    x"54",x"4F",x"52",x"45",x"8C",x"45",x"54",x"49", -- 0x3420
    x"52",x"51",x"8E",x"45",x"54",x"4E",x"4D",x"49", -- 0x3428
    x"8F",x"45",x"54",x"55",x"52",x"4E",x"90",x"49", -- 0x3430
    x"47",x"48",x"54",x"24",x"28",x"E3",x"4E",x"44", -- 0x3438
    x"28",x"C9",x"55",x"4E",x"8A",x"00",x"41",x"44", -- 0x3440
    x"44",x"28",x"D2",x"41",x"56",x"45",x"98",x"47", -- 0x3448
    x"4E",x"28",x"C2",x"49",x"4E",x"28",x"CD",x"50", -- 0x3450
    x"43",x"28",x"AE",x"51",x"52",x"28",x"C8",x"54", -- 0x3458
    x"45",x"50",x"B1",x"54",x"4F",x"50",x"92",x"54", -- 0x3460
    x"52",x"24",x"28",x"D4",x"57",x"41",x"50",x"A6", -- 0x3468
    x"00",x"41",x"42",x"28",x"AB",x"41",x"4E",x"28", -- 0x3470
    x"CE",x"48",x"45",x"4E",x"AF",x"4F",x"AC",x"57", -- 0x3478
    x"4F",x"50",x"49",x"E0",x"00",x"43",x"41",x"53", -- 0x3480
    x"45",x"24",x"28",x"D7",x"4E",x"54",x"49",x"4C", -- 0x3488
    x"B2",x"53",x"52",x"28",x"C5",x"00",x"41",x"4C", -- 0x3490
    x"28",x"D5",x"41",x"52",x"50",x"54",x"52",x"28", -- 0x3498
    x"E1",x"00",x"41",x"49",x"54",x"96",x"48",x"49", -- 0x34A0
    x"4C",x"45",x"B3",x"49",x"44",x"54",x"48",x"A4", -- 0x34A8
    x"00",x"B9",x"00",x"03",x"45",x"7B",x"F3",x"03", -- 0x34B0
    x"46",x"88",x"F3",x"04",x"4E",x"EB",x"F3",x"04", -- 0x34B8
    x"44",x"62",x"F3",x"05",x"49",x"A8",x"F3",x"03", -- 0x34C0
    x"44",x"71",x"F3",x"04",x"52",x"17",x"F4",x"03", -- 0x34C8
    x"4C",x"C6",x"F3",x"03",x"44",x"66",x"F3",x"04", -- 0x34D0
    x"47",x"98",x"F3",x"03",x"52",x"42",x"F4",x"02", -- 0x34D8
    x"49",x"A3",x"F3",x"07",x"52",x"1E",x"F4",x"05", -- 0x34E0
    x"47",x"93",x"F3",x"06",x"52",x"25",x"F4",x"06", -- 0x34E8
    x"52",x"2B",x"F4",x"06",x"52",x"31",x"F4",x"03", -- 0x34F0
    x"52",x"1B",x"F4",x"04",x"53",x"63",x"F4",x"02", -- 0x34F8
    x"4F",x"FD",x"F3",x"04",x"4E",x"F5",x"F3",x"03", -- 0x3500
    x"49",x"A5",x"F3",x"04",x"57",x"A2",x"F4",x"04", -- 0x3508
    x"4C",x"CD",x"F3",x"04",x"53",x"4B",x"F4",x"03", -- 0x3510
    x"44",x"6E",x"F3",x"04",x"50",x"09",x"F4",x"04", -- 0x3518
    x"44",x"74",x"F3",x"04",x"43",x"4B",x"F3",x"02", -- 0x3520
    x"44",x"78",x"F3",x"04",x"4C",x"D5",x"F3",x"05", -- 0x3528
    x"50",x"11",x"F4",x"04",x"43",x"59",x"F3",x"04", -- 0x3530
    x"4C",x"C9",x"F3",x"05",x"43",x"54",x"F3",x"03", -- 0x3538
    x"4E",x"E8",x"F3",x"05",x"57",x"AB",x"F4",x"03", -- 0x3540
    x"47",x"90",x"F3",x"04",x"53",x"6C",x"F4",x"06", -- 0x3548
    x"42",x"3D",x"F3",x"06",x"42",x"37",x"F3",x"03", -- 0x3550
    x"49",x"B1",x"F3",x"03",x"4E",x"EF",x"F3",x"04", -- 0x3558
    x"54",x"71",x"F4",x"02",x"54",x"7D",x"F4",x"02", -- 0x3560
    x"46",x"86",x"F3",x"04",x"53",x"57",x"F4",x"04", -- 0x3568
    x"54",x"79",x"F4",x"03",x"4E",x"F2",x"F3",x"04", -- 0x3570
    x"53",x"5F",x"F4",x"05",x"55",x"8C",x"F4",x"05", -- 0x3578
    x"57",x"A6",x"F4",x"03",x"4F",x"FA",x"F3",x"01", -- 0x3580
    x"2B",x"00",x"00",x"01",x"2D",x"00",x"00",x"01", -- 0x3588
    x"2A",x"00",x"00",x"01",x"2F",x"00",x"00",x"01", -- 0x3590
    x"5E",x"00",x"00",x"03",x"41",x"26",x"F3",x"03", -- 0x3598
    x"45",x"7E",x"F3",x"02",x"4F",x"FF",x"F3",x"02", -- 0x35A0
    x"3E",x"1C",x"F3",x"02",x"3C",x"16",x"F3",x"01", -- 0x35A8
    x"3E",x"00",x"00",x"01",x"3D",x"00",x"00",x"01", -- 0x35B0
    x"3C",x"00",x"00",x"04",x"53",x"4F",x"F4",x"04", -- 0x35B8
    x"49",x"AD",x"F3",x"04",x"41",x"22",x"F3",x"04", -- 0x35C0
    x"55",x"91",x"F4",x"04",x"46",x"8B",x"F3",x"04", -- 0x35C8
    x"50",x"0D",x"F4",x"04",x"53",x"5B",x"F4",x"04", -- 0x35D0
    x"52",x"3E",x"F4",x"04",x"4C",x"D1",x"F3",x"04", -- 0x35D8
    x"45",x"81",x"F3",x"04",x"43",x"5D",x"F3",x"04", -- 0x35E0
    x"53",x"53",x"F4",x"04",x"54",x"75",x"F4",x"04", -- 0x35E8
    x"41",x"2D",x"F3",x"05",x"50",x"02",x"F4",x"05", -- 0x35F0
    x"44",x"69",x"F3",x"05",x"53",x"46",x"F4",x"04", -- 0x35F8
    x"4C",x"C2",x"F3",x"05",x"53",x"67",x"F4",x"04", -- 0x3600
    x"56",x"96",x"F4",x"04",x"41",x"29",x"F3",x"07", -- 0x3608
    x"55",x"85",x"F4",x"07",x"4C",x"B5",x"F3",x"05", -- 0x3610
    x"43",x"4F",x"F3",x"05",x"48",x"9D",x"F3",x"05", -- 0x3618
    x"42",x"32",x"F3",x"07",x"42",x"43",x"F3",x"04", -- 0x3620
    x"4D",x"DA",x"F3",x"04",x"4D",x"E3",x"F3",x"02", -- 0x3628
    x"50",x"07",x"F4",x"05",x"54",x"7F",x"F4",x"07", -- 0x3630
    x"56",x"9A",x"F4",x"06",x"4C",x"BC",x"F3",x"07", -- 0x3638
    x"52",x"37",x"F4",x"05",x"4D",x"DE",x"F3",x"6B", -- 0x3640
    x"F6",x"7C",x"F6",x"83",x"F6",x"98",x"F6",x"A4", -- 0x3648
    x"F6",x"B2",x"F6",x"BB",x"F6",x"C9",x"F6",x"DD", -- 0x3650
    x"F6",x"EA",x"F6",x"FB",x"F6",x"0A",x"F7",x"19", -- 0x3658
    x"F7",x"27",x"F7",x"37",x"F7",x"4A",x"F7",x"59", -- 0x3660
    x"F7",x"6C",x"F7",x"4E",x"45",x"58",x"54",x"20", -- 0x3668
    x"77",x"69",x"74",x"68",x"6F",x"75",x"74",x"20", -- 0x3670
    x"46",x"4F",x"52",x"00",x"53",x"79",x"6E",x"74", -- 0x3678
    x"61",x"78",x"00",x"52",x"45",x"54",x"55",x"52", -- 0x3680
    x"4E",x"20",x"77",x"69",x"74",x"68",x"6F",x"75", -- 0x3688
    x"74",x"20",x"47",x"4F",x"53",x"55",x"42",x"00", -- 0x3690
    x"4F",x"75",x"74",x"20",x"6F",x"66",x"20",x"44", -- 0x3698
    x"41",x"54",x"41",x"00",x"46",x"75",x"6E",x"63", -- 0x36A0
    x"74",x"69",x"6F",x"6E",x"20",x"63",x"61",x"6C", -- 0x36A8
    x"6C",x"00",x"4F",x"76",x"65",x"72",x"66",x"6C", -- 0x36B0
    x"6F",x"77",x"00",x"4F",x"75",x"74",x"20",x"6F", -- 0x36B8
    x"66",x"20",x"6D",x"65",x"6D",x"6F",x"72",x"79", -- 0x36C0
    x"00",x"55",x"6E",x"64",x"65",x"66",x"69",x"6E", -- 0x36C8
    x"65",x"64",x"20",x"73",x"74",x"61",x"74",x"65", -- 0x36D0
    x"6D",x"65",x"6E",x"74",x"00",x"41",x"72",x"72", -- 0x36D8
    x"61",x"79",x"20",x"62",x"6F",x"75",x"6E",x"64", -- 0x36E0
    x"73",x"00",x"44",x"6F",x"75",x"62",x"6C",x"65", -- 0x36E8
    x"20",x"64",x"69",x"6D",x"65",x"6E",x"73",x"69", -- 0x36F0
    x"6F",x"6E",x"00",x"44",x"69",x"76",x"69",x"64", -- 0x36F8
    x"65",x"20",x"62",x"79",x"20",x"7A",x"65",x"72", -- 0x3700
    x"6F",x"00",x"49",x"6C",x"6C",x"65",x"67",x"61", -- 0x3708
    x"6C",x"20",x"64",x"69",x"72",x"65",x"63",x"74", -- 0x3710
    x"00",x"54",x"79",x"70",x"65",x"20",x"6D",x"69", -- 0x3718
    x"73",x"6D",x"61",x"74",x"63",x"68",x"00",x"53", -- 0x3720
    x"74",x"72",x"69",x"6E",x"67",x"20",x"74",x"6F", -- 0x3728
    x"6F",x"20",x"6C",x"6F",x"6E",x"67",x"00",x"53", -- 0x3730
    x"74",x"72",x"69",x"6E",x"67",x"20",x"74",x"6F", -- 0x3738
    x"6F",x"20",x"63",x"6F",x"6D",x"70",x"6C",x"65", -- 0x3740
    x"78",x"00",x"43",x"61",x"6E",x"27",x"74",x"20", -- 0x3748
    x"63",x"6F",x"6E",x"74",x"69",x"6E",x"75",x"65", -- 0x3750
    x"00",x"55",x"6E",x"64",x"65",x"66",x"69",x"6E", -- 0x3758
    x"65",x"64",x"20",x"66",x"75",x"6E",x"63",x"74", -- 0x3760
    x"69",x"6F",x"6E",x"00",x"4C",x"4F",x"4F",x"50", -- 0x3768
    x"20",x"77",x"69",x"74",x"68",x"6F",x"75",x"74", -- 0x3770
    x"20",x"44",x"4F",x"00",x"0D",x"0A",x"42",x"72", -- 0x3778
    x"65",x"61",x"6B",x"00",x"20",x"45",x"72",x"72", -- 0x3780
    x"6F",x"72",x"00",x"20",x"69",x"6E",x"20",x"6C", -- 0x3788
    x"69",x"6E",x"65",x"20",x"00",x"0D",x"0A",x"52", -- 0x3790
    x"65",x"61",x"64",x"79",x"0D",x"0A",x"00",x"20", -- 0x3798
    x"45",x"78",x"74",x"72",x"61",x"20",x"69",x"67", -- 0x37A0
    x"6E",x"6F",x"72",x"65",x"64",x"0D",x"0A",x"00", -- 0x37A8
    x"20",x"52",x"65",x"64",x"6F",x"20",x"66",x"72", -- 0x37B0
    x"6F",x"6D",x"20",x"73",x"74",x"61",x"72",x"74", -- 0x37B8
    x"0D",x"0A",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
    x"5A",x"4D",x"32",x"3A",x"20",x"53",x"74",x"61", -- 0x3800
    x"72",x"74",x"69",x"6E",x"67",x"2E",x"2E",x"2E", -- 0x3808
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3810
    x"00",x"00",x"00",x"00",x"00",x"09",x"60",x"00", -- 0x3818
    x"00",x"00",x"00",x"00",x"00",x"51",x"31",x"00", -- 0x3820
    x"00",x"00",x"5A",x"53",x"41",x"57",x"32",x"00", -- 0x3828
    x"00",x"43",x"58",x"44",x"45",x"34",x"33",x"00", -- 0x3830
    x"00",x"20",x"56",x"46",x"54",x"52",x"35",x"00", -- 0x3838
    x"00",x"4E",x"42",x"48",x"47",x"59",x"36",x"00", -- 0x3840
    x"00",x"00",x"4D",x"4A",x"55",x"37",x"38",x"00", -- 0x3848
    x"00",x"2C",x"4B",x"49",x"4F",x"30",x"39",x"00", -- 0x3850
    x"00",x"2E",x"2F",x"4C",x"3B",x"50",x"2D",x"00", -- 0x3858
    x"00",x"00",x"00",x"00",x"5B",x"3D",x"00",x"00", -- 0x3860
    x"00",x"00",x"0D",x"5D",x"00",x"5C",x"00",x"00", -- 0x3868
    x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x3870
    x"00",x"31",x"00",x"34",x"37",x"00",x"00",x"00", -- 0x3878
    x"30",x"2E",x"32",x"35",x"36",x"38",x"03",x"00", -- 0x3880
    x"00",x"2B",x"33",x"2D",x"2A",x"39",x"00",x"00", -- 0x3888
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3890
    x"00",x"00",x"00",x"00",x"00",x"09",x"AC",x"00", -- 0x3898
    x"00",x"00",x"00",x"00",x"00",x"71",x"21",x"00", -- 0x38A0
    x"00",x"00",x"7A",x"73",x"61",x"77",x"22",x"00", -- 0x38A8
    x"00",x"63",x"78",x"64",x"65",x"24",x"A3",x"00", -- 0x38B0
    x"00",x"20",x"76",x"66",x"74",x"72",x"25",x"00", -- 0x38B8
    x"00",x"6E",x"62",x"68",x"67",x"79",x"5E",x"00", -- 0x38C0
    x"00",x"00",x"6D",x"6A",x"75",x"26",x"2A",x"00", -- 0x38C8
    x"00",x"3C",x"6B",x"69",x"6F",x"29",x"28",x"00", -- 0x38D0
    x"00",x"3E",x"3F",x"6C",x"3A",x"70",x"5F",x"00", -- 0x38D8
    x"00",x"00",x"00",x"00",x"5B",x"2B",x"00",x"00", -- 0x38E0
    x"00",x"00",x"0D",x"5D",x"00",x"5C",x"00",x"00", -- 0x38E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x38F0
    x"00",x"31",x"00",x"34",x"37",x"00",x"00",x"00", -- 0x38F8
    x"30",x"2E",x"32",x"35",x"36",x"38",x"03",x"00", -- 0x3900
    x"00",x"2B",x"33",x"2D",x"2A",x"39",x"00",x"00", -- 0x3908
    x"D8",x"A2",x"FF",x"9A",x"20",x"34",x"F9",x"A9", -- 0x3910
    x"00",x"85",x"E8",x"A2",x"10",x"BD",x"FF",x"F7", -- 0x3918
    x"9D",x"FF",x"BF",x"CA",x"D0",x"F7",x"A0",x"08", -- 0x3920
    x"B9",x"C2",x"FA",x"99",x"04",x"02",x"88",x"D0", -- 0x3928
    x"F7",x"4C",x"00",x"D0",x"A9",x"C0",x"85",x"EE", -- 0x3930
    x"A9",x"00",x"85",x"ED",x"A8",x"A2",x"09",x"91", -- 0x3938
    x"ED",x"C8",x"D0",x"FB",x"E6",x"EE",x"CA",x"D0", -- 0x3940
    x"F6",x"A2",x"60",x"91",x"ED",x"C8",x"CA",x"D0", -- 0x3948
    x"FA",x"A9",x"C0",x"85",x"EE",x"A9",x"00",x"85", -- 0x3950
    x"ED",x"85",x"EA",x"85",x"E9",x"60",x"A9",x"C0", -- 0x3958
    x"85",x"EE",x"85",x"EC",x"A9",x"50",x"85",x"EB", -- 0x3960
    x"A9",x"00",x"85",x"ED",x"A8",x"A2",x"09",x"B1", -- 0x3968
    x"EB",x"91",x"ED",x"C8",x"D0",x"F9",x"E6",x"EC", -- 0x3970
    x"E6",x"EE",x"CA",x"D0",x"F2",x"A2",x"10",x"B1", -- 0x3978
    x"EB",x"91",x"ED",x"C8",x"CA",x"D0",x"F8",x"A5", -- 0x3980
    x"ED",x"69",x"0F",x"85",x"ED",x"A2",x"50",x"A9", -- 0x3988
    x"00",x"A8",x"91",x"ED",x"C8",x"CA",x"D0",x"FA", -- 0x3990
    x"C6",x"E9",x"60",x"85",x"E5",x"8A",x"48",x"98", -- 0x3998
    x"48",x"A5",x"E5",x"C9",x"0A",x"F0",x"28",x"C9", -- 0x39A0
    x"0D",x"F0",x"34",x"C9",x"08",x"F0",x"42",x"A0", -- 0x39A8
    x"00",x"91",x"ED",x"18",x"A5",x"ED",x"69",x"01", -- 0x39B0
    x"85",x"ED",x"90",x"02",x"E6",x"EE",x"A5",x"EA", -- 0x39B8
    x"E6",x"EA",x"C9",x"50",x"90",x"06",x"A9",x"00", -- 0x39C0
    x"85",x"EA",x"E6",x"E9",x"4C",x"07",x"FA",x"18", -- 0x39C8
    x"A5",x"ED",x"69",x"50",x"85",x"ED",x"90",x"02", -- 0x39D0
    x"E6",x"EE",x"E6",x"E9",x"4C",x"07",x"FA",x"38", -- 0x39D8
    x"A5",x"ED",x"E5",x"EA",x"85",x"ED",x"B0",x"02", -- 0x39E0
    x"C6",x"EE",x"A9",x"00",x"85",x"EA",x"4C",x"07", -- 0x39E8
    x"FA",x"A5",x"EA",x"F0",x"12",x"C6",x"EA",x"38", -- 0x39F0
    x"A5",x"ED",x"E9",x"01",x"85",x"ED",x"B0",x"02", -- 0x39F8
    x"C6",x"EE",x"A9",x"00",x"A8",x"91",x"ED",x"A5", -- 0x3A00
    x"E9",x"C9",x"1E",x"D0",x"03",x"20",x"5E",x"F9", -- 0x3A08
    x"A5",x"EA",x"8D",x"FC",x"CB",x"A5",x"E9",x"8D", -- 0x3A10
    x"FD",x"CB",x"68",x"A8",x"68",x"AA",x"A5",x"E5", -- 0x3A18
    x"60",x"85",x"E5",x"8A",x"48",x"A5",x"E5",x"A5", -- 0x3A20
    x"E7",x"85",x"E5",x"F0",x"08",x"A2",x"00",x"86", -- 0x3A28
    x"E7",x"38",x"4C",x"36",x"FA",x"18",x"68",x"AA", -- 0x3A30
    x"A5",x"E5",x"60",x"48",x"8A",x"48",x"AD",x"00", -- 0x3A38
    x"CC",x"AA",x"C9",x"F0",x"F0",x"67",x"C9",x"80", -- 0x3A40
    x"F0",x"6C",x"A9",x"02",x"24",x"E8",x"D0",x"26", -- 0x3A48
    x"A9",x"01",x"24",x"E8",x"D0",x"4E",x"E0",x"12", -- 0x3A50
    x"F0",x"38",x"E0",x"59",x"F0",x"34",x"A9",x"10", -- 0x3A58
    x"24",x"E8",x"D0",x"0A",x"BD",x"10",x"F8",x"85", -- 0x3A60
    x"E7",x"85",x"E6",x"4C",x"BF",x"FA",x"BD",x"90", -- 0x3A68
    x"F8",x"85",x"E7",x"4C",x"BF",x"FA",x"A5",x"E8", -- 0x3A70
    x"29",x"FD",x"85",x"E8",x"E0",x"12",x"F0",x"1B", -- 0x3A78
    x"E0",x"59",x"F0",x"17",x"BD",x"10",x"F8",x"C5", -- 0x3A80
    x"E6",x"D0",x"34",x"A9",x"00",x"85",x"E6",x"4C", -- 0x3A88
    x"BF",x"FA",x"A5",x"E8",x"09",x"10",x"85",x"E8", -- 0x3A90
    x"4C",x"BF",x"FA",x"A5",x"E8",x"29",x"EF",x"85", -- 0x3A98
    x"E8",x"4C",x"BF",x"FA",x"A5",x"E8",x"29",x"FE", -- 0x3AA0
    x"85",x"E8",x"4C",x"BF",x"FA",x"A5",x"E8",x"09", -- 0x3AA8
    x"02",x"85",x"E8",x"4C",x"BF",x"FA",x"A5",x"E8", -- 0x3AB0
    x"09",x"01",x"85",x"E8",x"4C",x"BF",x"FA",x"68", -- 0x3AB8
    x"AA",x"68",x"40",x"21",x"FA",x"9B",x"F9",x"3A", -- 0x3AC0
    x"FA",x"3A",x"FA",x"00",x"00",x"00",x"00",x"00", -- 0x3AC8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF8
    x"20",x"34",x"F9",x"A0",x"00",x"A9",x"DA",x"91", -- 0x3B00
    x"ED",x"E6",x"ED",x"A9",x"C4",x"A0",x"4E",x"20", -- 0x3B08
    x"46",x"FF",x"A9",x"BF",x"91",x"ED",x"E6",x"ED", -- 0x3B10
    x"A9",x"B3",x"A0",x"1C",x"20",x"5B",x"FF",x"A9", -- 0x3B18
    x"C0",x"91",x"ED",x"E6",x"ED",x"A9",x"C4",x"A0", -- 0x3B20
    x"4E",x"20",x"46",x"FF",x"A9",x"D9",x"91",x"ED", -- 0x3B28
    x"A9",x"9F",x"85",x"ED",x"A9",x"C0",x"85",x"EE", -- 0x3B30
    x"A9",x"B3",x"A0",x"1C",x"20",x"5B",x"FF",x"A9", -- 0x3B38
    x"C4",x"85",x"EC",x"85",x"EE",x"A9",x"CE",x"85", -- 0x3B40
    x"EB",x"85",x"ED",x"A9",x"01",x"8D",x"FC",x"FB", -- 0x3B48
    x"8D",x"FD",x"FB",x"A0",x"0A",x"A9",x"CD",x"20", -- 0x3B50
    x"46",x"FF",x"A5",x"E6",x"C9",x"57",x"F0",x"11", -- 0x3B58
    x"C9",x"41",x"F0",x"12",x"C9",x"53",x"F0",x"13", -- 0x3B60
    x"C9",x"44",x"D0",x"14",x"A9",x"01",x"4C",x"7D", -- 0x3B68
    x"FB",x"A9",x"00",x"4C",x"7D",x"FB",x"A9",x"03", -- 0x3B70
    x"4C",x"7D",x"FB",x"A9",x"02",x"8D",x"FE",x"FB", -- 0x3B78
    x"A0",x"00",x"B1",x"ED",x"F0",x"03",x"4C",x"00", -- 0x3B80
    x"FB",x"AD",x"FD",x"FB",x"18",x"2A",x"2A",x"6D", -- 0x3B88
    x"FE",x"FB",x"AA",x"BD",x"E8",x"FB",x"F0",x"C2", -- 0x3B90
    x"91",x"ED",x"AE",x"FE",x"FB",x"8E",x"FD",x"FB", -- 0x3B98
    x"BD",x"F8",x"FB",x"10",x"02",x"A0",x"FF",x"65", -- 0x3BA0
    x"ED",x"85",x"ED",x"98",x"65",x"EE",x"85",x"EE", -- 0x3BA8
    x"AD",x"FC",x"FB",x"18",x"2A",x"2A",x"AA",x"A0", -- 0x3BB0
    x"00",x"B1",x"EB",x"CA",x"88",x"E8",x"C8",x"DD", -- 0x3BB8
    x"E8",x"FB",x"D0",x"F9",x"8C",x"FC",x"FB",x"BE", -- 0x3BC0
    x"F8",x"FB",x"A9",x"00",x"A8",x"91",x"EB",x"E0", -- 0x3BC8
    x"80",x"90",x"02",x"A0",x"FF",x"8A",x"18",x"65", -- 0x3BD0
    x"EB",x"85",x"EB",x"98",x"65",x"EC",x"85",x"EC", -- 0x3BD8
    x"A9",x"FF",x"20",x"76",x"FF",x"4C",x"5A",x"FB", -- 0x3BE0
    x"BA",x"C9",x"00",x"BB",x"BC",x"CD",x"BB",x"00", -- 0x3BE8
    x"00",x"C8",x"BA",x"BC",x"C8",x"00",x"C9",x"CD", -- 0x3BF0
    x"B0",x"01",x"50",x"FF",x"01",x"01",x"01",x"00", -- 0x3BF8
    x"A9",x"C0",x"8D",x"09",x"10",x"20",x"08",x"FE", -- 0x3C00
    x"20",x"DB",x"FE",x"20",x"A7",x"FD",x"A2",x"14", -- 0x3C08
    x"20",x"11",x"FD",x"AD",x"09",x"10",x"20",x"76", -- 0x3C10
    x"FF",x"A5",x"E6",x"C9",x"03",x"D0",x"03",x"4C", -- 0x3C18
    x"08",x"FD",x"C9",x"41",x"D0",x"09",x"CE",x"02", -- 0x3C20
    x"10",x"EE",x"0D",x"10",x"4C",x"39",x"FC",x"C9", -- 0x3C28
    x"44",x"D0",x"06",x"EE",x"02",x"10",x"EE",x"0E", -- 0x3C30
    x"10",x"AD",x"02",x"10",x"C9",x"01",x"B0",x"05", -- 0x3C38
    x"A9",x"01",x"8D",x"02",x"10",x"C9",x"45",x"90", -- 0x3C40
    x"05",x"A9",x"45",x"8D",x"02",x"10",x"CD",x"03", -- 0x3C48
    x"10",x"F0",x"09",x"20",x"A7",x"FD",x"AD",x"02", -- 0x3C50
    x"10",x"8D",x"03",x"10",x"EE",x"06",x"10",x"AD", -- 0x3C58
    x"06",x"10",x"29",x"01",x"F0",x"AD",x"A9",x"00", -- 0x3C60
    x"A8",x"91",x"ED",x"AD",x"00",x"10",x"20",x"27", -- 0x3C68
    x"FD",x"8D",x"00",x"10",x"AD",x"01",x"10",x"20", -- 0x3C70
    x"27",x"FD",x"8D",x"01",x"10",x"38",x"A5",x"ED", -- 0x3C78
    x"E9",x"C0",x"A5",x"EE",x"E9",x"C8",x"90",x"13", -- 0x3C80
    x"A9",x"00",x"AE",x"0A",x"10",x"9D",x"9A",x"C0", -- 0x3C88
    x"CA",x"8E",x"0A",x"10",x"F0",x"3C",x"A2",x"0A", -- 0x3C90
    x"20",x"11",x"FD",x"A0",x"00",x"B1",x"ED",x"F0", -- 0x3C98
    x"20",x"20",x"72",x"FD",x"D0",x"03",x"20",x"C4", -- 0x3CA0
    x"FD",x"38",x"A9",x"00",x"ED",x"00",x"10",x"8D", -- 0x3CA8
    x"00",x"10",x"20",x"27",x"FD",x"38",x"A9",x"00", -- 0x3CB0
    x"ED",x"01",x"10",x"8D",x"01",x"10",x"20",x"27", -- 0x3CB8
    x"FD",x"A9",x"02",x"A0",x"00",x"91",x"ED",x"AD", -- 0x3CC0
    x"08",x"10",x"D0",x"03",x"4C",x"08",x"FC",x"4C", -- 0x3CC8
    x"13",x"FC",x"A9",x"B4",x"85",x"EB",x"A9",x"FF", -- 0x3CD0
    x"85",x"EC",x"A9",x"FE",x"85",x"ED",x"A9",x"C1", -- 0x3CD8
    x"85",x"EE",x"20",x"89",x"FF",x"18",x"A5",x"ED", -- 0x3CE0
    x"69",x"4C",x"85",x"ED",x"90",x"02",x"E6",x"EE", -- 0x3CE8
    x"A9",x"C7",x"85",x"EB",x"A9",x"FF",x"85",x"EC", -- 0x3CF0
    x"20",x"89",x"FF",x"A5",x"E6",x"C9",x"03",x"F0", -- 0x3CF8
    x"07",x"C9",x"0D",x"D0",x"CD",x"4C",x"00",x"FC", -- 0x3D00
    x"20",x"34",x"F9",x"A9",x"FF",x"8D",x"FE",x"CB", -- 0x3D08
    x"60",x"A9",x"00",x"A8",x"91",x"ED",x"A9",x"FF", -- 0x3D10
    x"20",x"76",x"FF",x"A9",x"02",x"91",x"ED",x"A9", -- 0x3D18
    x"FF",x"20",x"76",x"FF",x"CA",x"D0",x"EA",x"8D", -- 0x3D20
    x"0B",x"10",x"C9",x"80",x"B0",x"08",x"A9",x"00", -- 0x3D28
    x"8D",x"0C",x"10",x"4C",x"3B",x"FD",x"A9",x"FF", -- 0x3D30
    x"8D",x"0C",x"10",x"18",x"A5",x"ED",x"6D",x"0B", -- 0x3D38
    x"10",x"85",x"ED",x"A5",x"EE",x"6D",x"0C",x"10", -- 0x3D40
    x"85",x"EE",x"A0",x"00",x"B1",x"ED",x"D0",x"04", -- 0x3D48
    x"AD",x"0B",x"10",x"60",x"20",x"72",x"FD",x"D0", -- 0x3D50
    x"03",x"20",x"C4",x"FD",x"38",x"A5",x"ED",x"ED", -- 0x3D58
    x"0B",x"10",x"85",x"ED",x"A5",x"EE",x"ED",x"0C", -- 0x3D60
    x"10",x"85",x"EE",x"38",x"A9",x"00",x"ED",x"0B", -- 0x3D68
    x"10",x"60",x"A5",x"ED",x"8D",x"07",x"10",x"29", -- 0x3D70
    x"FC",x"85",x"ED",x"A2",x"00",x"A0",x"04",x"88", -- 0x3D78
    x"B1",x"ED",x"C9",x"DB",x"F0",x"0F",x"C9",x"B0", -- 0x3D80
    x"F0",x"0B",x"C9",x"B1",x"F0",x"07",x"C9",x"B2", -- 0x3D88
    x"F0",x"03",x"4C",x"9B",x"FD",x"A2",x"01",x"A9", -- 0x3D90
    x"00",x"91",x"ED",x"C0",x"00",x"D0",x"E0",x"AD", -- 0x3D98
    x"07",x"10",x"85",x"ED",x"E0",x"01",x"60",x"AE", -- 0x3DA0
    x"03",x"10",x"A0",x"0A",x"A9",x"00",x"9D",x"C0", -- 0x3DA8
    x"C8",x"E8",x"88",x"D0",x"F9",x"AE",x"02",x"10", -- 0x3DB0
    x"A0",x"0A",x"A9",x"CD",x"9D",x"C0",x"C8",x"E8", -- 0x3DB8
    x"88",x"D0",x"F9",x"60",x"CE",x"08",x"10",x"18", -- 0x3DC0
    x"AD",x"5C",x"C0",x"69",x"05",x"C9",x"3A",x"B0", -- 0x3DC8
    x"04",x"8D",x"5C",x"C0",x"60",x"38",x"E9",x"0A", -- 0x3DD0
    x"8D",x"5C",x"C0",x"CE",x"09",x"10",x"18",x"AD", -- 0x3DD8
    x"5B",x"C0",x"69",x"01",x"C9",x"3A",x"B0",x"04", -- 0x3DE0
    x"8D",x"5B",x"C0",x"60",x"A9",x"30",x"8D",x"5B", -- 0x3DE8
    x"C0",x"18",x"AD",x"5A",x"C0",x"69",x"01",x"C9", -- 0x3DF0
    x"3A",x"B0",x"04",x"8D",x"5A",x"C0",x"60",x"A9", -- 0x3DF8
    x"30",x"8D",x"5A",x"C0",x"EE",x"59",x"C0",x"60", -- 0x3E00
    x"20",x"34",x"F9",x"A9",x"00",x"8D",x"FE",x"CB", -- 0x3E08
    x"A8",x"A9",x"DA",x"91",x"ED",x"E6",x"ED",x"A9", -- 0x3E10
    x"C4",x"A0",x"4E",x"20",x"46",x"FF",x"A9",x"BF", -- 0x3E18
    x"91",x"ED",x"E6",x"ED",x"A9",x"B3",x"91",x"ED", -- 0x3E20
    x"E6",x"ED",x"E6",x"ED",x"A9",x"96",x"85",x"EB", -- 0x3E28
    x"A9",x"FF",x"85",x"EC",x"20",x"89",x"FF",x"A9", -- 0x3E30
    x"30",x"8D",x"5C",x"C0",x"8D",x"5B",x"C0",x"8D", -- 0x3E38
    x"5A",x"C0",x"8D",x"59",x"C0",x"18",x"A5",x"ED", -- 0x3E40
    x"69",x"1E",x"85",x"ED",x"A9",x"A4",x"85",x"EB", -- 0x3E48
    x"A9",x"FF",x"85",x"EC",x"20",x"89",x"FF",x"A5", -- 0x3E50
    x"ED",x"69",x"24",x"85",x"ED",x"A9",x"9D",x"85", -- 0x3E58
    x"EB",x"A9",x"FF",x"85",x"EC",x"20",x"89",x"FF", -- 0x3E60
    x"A0",x"00",x"A5",x"ED",x"69",x"07",x"85",x"ED", -- 0x3E68
    x"A9",x"02",x"91",x"ED",x"E6",x"ED",x"91",x"ED", -- 0x3E70
    x"E6",x"ED",x"91",x"ED",x"E6",x"ED",x"E6",x"ED", -- 0x3E78
    x"A9",x"B3",x"91",x"ED",x"E6",x"ED",x"A9",x"C3", -- 0x3E80
    x"91",x"ED",x"E6",x"ED",x"A9",x"C4",x"A0",x"4E", -- 0x3E88
    x"20",x"46",x"FF",x"A9",x"B4",x"91",x"ED",x"E6", -- 0x3E90
    x"ED",x"A9",x"B3",x"A0",x"1A",x"20",x"5B",x"FF", -- 0x3E98
    x"A9",x"3F",x"85",x"ED",x"A9",x"C1",x"85",x"EE", -- 0x3EA0
    x"A9",x"B3",x"A0",x"1A",x"20",x"5B",x"FF",x"A9", -- 0x3EA8
    x"10",x"85",x"ED",x"A9",x"C9",x"85",x"EE",x"A9", -- 0x3EB0
    x"C0",x"91",x"ED",x"E6",x"ED",x"A9",x"C4",x"A0", -- 0x3EB8
    x"4E",x"20",x"46",x"FF",x"A9",x"D9",x"91",x"ED", -- 0x3EC0
    x"A9",x"D7",x"85",x"ED",x"A9",x"C4",x"85",x"EE", -- 0x3EC8
    x"A9",x"01",x"8D",x"03",x"10",x"A9",x"03",x"8D", -- 0x3ED0
    x"0A",x"10",x"60",x"A9",x"00",x"A8",x"91",x"ED", -- 0x3ED8
    x"A9",x"91",x"85",x"ED",x"A9",x"C1",x"85",x"EE", -- 0x3EE0
    x"A9",x"DB",x"A0",x"4E",x"20",x"46",x"FF",x"A9", -- 0x3EE8
    x"E1",x"85",x"ED",x"A9",x"C1",x"85",x"EE",x"A9", -- 0x3EF0
    x"B2",x"A0",x"4E",x"20",x"46",x"FF",x"A9",x"31", -- 0x3EF8
    x"85",x"ED",x"A9",x"C2",x"85",x"EE",x"A9",x"B1", -- 0x3F00
    x"A0",x"4E",x"20",x"46",x"FF",x"A9",x"81",x"85", -- 0x3F08
    x"ED",x"A9",x"C2",x"85",x"EE",x"A9",x"B0",x"A0", -- 0x3F10
    x"4E",x"20",x"46",x"FF",x"AD",x"0E",x"10",x"29", -- 0x3F18
    x"01",x"D0",x"02",x"A9",x"FF",x"8D",x"00",x"10", -- 0x3F20
    x"A9",x"B0",x"8D",x"01",x"10",x"AD",x"0D",x"10", -- 0x3F28
    x"29",x"07",x"38",x"69",x"D4",x"85",x"ED",x"A9", -- 0x3F30
    x"C4",x"85",x"EE",x"A9",x"50",x"8D",x"08",x"10", -- 0x3F38
    x"A9",x"25",x"8D",x"02",x"10",x"60",x"8C",x"07", -- 0x3F40
    x"10",x"88",x"91",x"ED",x"D0",x"FB",x"18",x"A5", -- 0x3F48
    x"ED",x"6D",x"07",x"10",x"85",x"ED",x"90",x"02", -- 0x3F50
    x"E6",x"EE",x"60",x"8D",x"07",x"10",x"98",x"AA", -- 0x3F58
    x"A0",x"00",x"AD",x"07",x"10",x"91",x"ED",x"18", -- 0x3F60
    x"A5",x"ED",x"69",x"50",x"85",x"ED",x"90",x"02", -- 0x3F68
    x"E6",x"EE",x"CA",x"D0",x"ED",x"60",x"8D",x"05", -- 0x3F70
    x"10",x"A9",x"00",x"8D",x"04",x"10",x"CE",x"04", -- 0x3F78
    x"10",x"D0",x"FB",x"CE",x"05",x"10",x"D0",x"F6", -- 0x3F80
    x"60",x"A0",x"00",x"B1",x"EB",x"F0",x"06",x"91", -- 0x3F88
    x"ED",x"C8",x"4C",x"8B",x"FF",x"60",x"53",x"63", -- 0x3F90
    x"6F",x"72",x"65",x"3A",x"00",x"4C",x"69",x"76", -- 0x3F98
    x"65",x"73",x"3A",x"00",x"42",x"20",x"52",x"20", -- 0x3FA0
    x"45",x"20",x"41",x"20",x"4B",x"20",x"4F",x"20", -- 0x3FA8
    x"55",x"20",x"54",x"00",x"20",x"47",x"20",x"41", -- 0x3FB0
    x"20",x"4D",x"20",x"45",x"20",x"20",x"4F",x"20", -- 0x3FB8
    x"56",x"20",x"45",x"20",x"52",x"20",x"00",x"20", -- 0x3FC0
    x"50",x"72",x"65",x"73",x"73",x"20",x"45",x"4E", -- 0x3FC8
    x"54",x"45",x"52",x"20",x"74",x"6F",x"20",x"74", -- 0x3FD0
    x"72",x"79",x"20",x"61",x"67",x"61",x"69",x"6E", -- 0x3FD8
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FF0
    x"00",x"00",x"10",x"F9",x"10",x"F9",x"3B",x"FA"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
