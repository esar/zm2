-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity character_rom is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of character_rom is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0000
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
    x"00",x"00",x"7E",x"81",x"A5",x"81",x"81",x"BD", -- 0x0010
    x"99",x"81",x"81",x"7E",x"00",x"00",x"00",x"00", -- 0x0018
    x"00",x"00",x"7E",x"FF",x"DB",x"FF",x"FF",x"C3", -- 0x0020
    x"E7",x"FF",x"FF",x"7E",x"00",x"00",x"00",x"00", -- 0x0028
    x"00",x"00",x"00",x"00",x"6C",x"FE",x"FE",x"FE", -- 0x0030
    x"FE",x"7C",x"38",x"10",x"00",x"00",x"00",x"00", -- 0x0038
    x"00",x"00",x"00",x"00",x"10",x"38",x"7C",x"FE", -- 0x0040
    x"7C",x"38",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x0048
    x"00",x"00",x"00",x"18",x"3C",x"3C",x"E7",x"E7", -- 0x0050
    x"E7",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"18",x"3C",x"7E",x"FF",x"FF", -- 0x0060
    x"7E",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3C", -- 0x0070
    x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0078
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"C3", -- 0x0080
    x"C3",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0088
    x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"42", -- 0x0090
    x"42",x"66",x"3C",x"00",x"00",x"00",x"00",x"00", -- 0x0098
    x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"99",x"BD", -- 0x00A0
    x"BD",x"99",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A8
    x"00",x"00",x"1E",x"0E",x"1A",x"32",x"78",x"CC", -- 0x00B0
    x"CC",x"CC",x"CC",x"78",x"00",x"00",x"00",x"00", -- 0x00B8
    x"00",x"00",x"3C",x"66",x"66",x"66",x"66",x"3C", -- 0x00C0
    x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x00C8
    x"00",x"00",x"3F",x"33",x"3F",x"30",x"30",x"30", -- 0x00D0
    x"30",x"70",x"F0",x"E0",x"00",x"00",x"00",x"00", -- 0x00D8
    x"00",x"00",x"7F",x"63",x"7F",x"63",x"63",x"63", -- 0x00E0
    x"63",x"67",x"E7",x"E6",x"C0",x"00",x"00",x"00", -- 0x00E8
    x"00",x"00",x"00",x"18",x"18",x"DB",x"3C",x"E7", -- 0x00F0
    x"3C",x"DB",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x00F8
    x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FE",x"F8", -- 0x0100
    x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00", -- 0x0108
    x"00",x"02",x"06",x"0E",x"1E",x"3E",x"FE",x"3E", -- 0x0110
    x"1E",x"0E",x"06",x"02",x"00",x"00",x"00",x"00", -- 0x0118
    x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18", -- 0x0120
    x"7E",x"3C",x"18",x"00",x"00",x"00",x"00",x"00", -- 0x0128
    x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"66", -- 0x0130
    x"66",x"00",x"66",x"66",x"00",x"00",x"00",x"00", -- 0x0138
    x"00",x"00",x"7F",x"DB",x"DB",x"DB",x"7B",x"1B", -- 0x0140
    x"1B",x"1B",x"1B",x"1B",x"00",x"00",x"00",x"00", -- 0x0148
    x"00",x"7C",x"C6",x"60",x"38",x"6C",x"C6",x"C6", -- 0x0150
    x"6C",x"38",x"0C",x"C6",x"7C",x"00",x"00",x"00", -- 0x0158
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0160
    x"FE",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"00", -- 0x0168
    x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18", -- 0x0170
    x"7E",x"3C",x"18",x"7E",x"00",x"00",x"00",x"00", -- 0x0178
    x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18", -- 0x0180
    x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x0188
    x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0190
    x"18",x"7E",x"3C",x"18",x"00",x"00",x"00",x"00", -- 0x0198
    x"00",x"00",x"00",x"00",x"00",x"18",x"0C",x"FE", -- 0x01A0
    x"0C",x"18",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01A8
    x"00",x"00",x"00",x"00",x"00",x"30",x"60",x"FE", -- 0x01B0
    x"60",x"30",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0", -- 0x01C0
    x"C0",x"FE",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01C8
    x"00",x"00",x"00",x"00",x"00",x"24",x"66",x"FF", -- 0x01D0
    x"66",x"24",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x01D8
    x"00",x"00",x"00",x"00",x"10",x"38",x"38",x"7C", -- 0x01E0
    x"7C",x"FE",x"FE",x"00",x"00",x"00",x"00",x"00", -- 0x01E8
    x"00",x"00",x"00",x"00",x"FE",x"FE",x"7C",x"7C", -- 0x01F0
    x"38",x"38",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x01F8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0200
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0208
    x"00",x"00",x"18",x"3C",x"3C",x"3C",x"18",x"18", -- 0x0210
    x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x0218
    x"00",x"66",x"66",x"66",x"24",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"6C",x"6C",x"FE",x"6C",x"6C", -- 0x0230
    x"6C",x"FE",x"6C",x"6C",x"00",x"00",x"00",x"00", -- 0x0238
    x"18",x"18",x"7C",x"C6",x"C2",x"C0",x"7C",x"06", -- 0x0240
    x"06",x"86",x"C6",x"7C",x"18",x"18",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"00",x"C2",x"C6",x"0C",x"18", -- 0x0250
    x"30",x"60",x"C6",x"86",x"00",x"00",x"00",x"00", -- 0x0258
    x"00",x"00",x"38",x"6C",x"6C",x"38",x"76",x"DC", -- 0x0260
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0268
    x"00",x"30",x"30",x"30",x"60",x"00",x"00",x"00", -- 0x0270
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0278
    x"00",x"00",x"0C",x"18",x"30",x"30",x"30",x"30", -- 0x0280
    x"30",x"30",x"18",x"0C",x"00",x"00",x"00",x"00", -- 0x0288
    x"00",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"0C", -- 0x0290
    x"0C",x"0C",x"18",x"30",x"00",x"00",x"00",x"00", -- 0x0298
    x"00",x"00",x"00",x"00",x"00",x"66",x"3C",x"FF", -- 0x02A0
    x"3C",x"66",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
    x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"7E", -- 0x02B0
    x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02C0
    x"00",x"18",x"18",x"18",x"30",x"00",x"00",x"00", -- 0x02C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E", -- 0x02D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02E0
    x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x02E8
    x"00",x"00",x"00",x"00",x"02",x"06",x"0C",x"18", -- 0x02F0
    x"30",x"60",x"C0",x"80",x"00",x"00",x"00",x"00", -- 0x02F8
    x"00",x"00",x"7C",x"C6",x"C6",x"CE",x"DE",x"F6", -- 0x0300
    x"E6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0308
    x"00",x"00",x"18",x"38",x"78",x"18",x"18",x"18", -- 0x0310
    x"18",x"18",x"18",x"7E",x"00",x"00",x"00",x"00", -- 0x0318
    x"00",x"00",x"7C",x"C6",x"06",x"0C",x"18",x"30", -- 0x0320
    x"60",x"C0",x"C6",x"FE",x"00",x"00",x"00",x"00", -- 0x0328
    x"00",x"00",x"7C",x"C6",x"06",x"06",x"3C",x"06", -- 0x0330
    x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0338
    x"00",x"00",x"0C",x"1C",x"3C",x"6C",x"CC",x"FE", -- 0x0340
    x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"00", -- 0x0348
    x"00",x"00",x"FE",x"C0",x"C0",x"C0",x"FC",x"06", -- 0x0350
    x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0358
    x"00",x"00",x"38",x"60",x"C0",x"C0",x"FC",x"C6", -- 0x0360
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0368
    x"00",x"00",x"FE",x"C6",x"06",x"06",x"0C",x"18", -- 0x0370
    x"30",x"30",x"30",x"30",x"00",x"00",x"00",x"00", -- 0x0378
    x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"7C",x"C6", -- 0x0380
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0388
    x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"7E",x"06", -- 0x0390
    x"06",x"06",x"0C",x"78",x"00",x"00",x"00",x"00", -- 0x0398
    x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00", -- 0x03A0
    x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
    x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00", -- 0x03B0
    x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00", -- 0x03B8
    x"00",x"00",x"00",x"06",x"0C",x"18",x"30",x"60", -- 0x03C0
    x"30",x"18",x"0C",x"06",x"00",x"00",x"00",x"00", -- 0x03C8
    x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00", -- 0x03D0
    x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
    x"00",x"00",x"00",x"60",x"30",x"18",x"0C",x"06", -- 0x03E0
    x"0C",x"18",x"30",x"60",x"00",x"00",x"00",x"00", -- 0x03E8
    x"00",x"00",x"7C",x"C6",x"C6",x"0C",x"18",x"18", -- 0x03F0
    x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x03F8
    x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"DE",x"DE", -- 0x0400
    x"DE",x"DC",x"C0",x"7C",x"00",x"00",x"00",x"00", -- 0x0408
    x"00",x"00",x"10",x"38",x"6C",x"C6",x"C6",x"FE", -- 0x0410
    x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x0418
    x"00",x"00",x"FC",x"66",x"66",x"66",x"7C",x"66", -- 0x0420
    x"66",x"66",x"66",x"FC",x"00",x"00",x"00",x"00", -- 0x0428
    x"00",x"00",x"3C",x"66",x"C2",x"C0",x"C0",x"C0", -- 0x0430
    x"C0",x"C2",x"66",x"3C",x"00",x"00",x"00",x"00", -- 0x0438
    x"00",x"00",x"F8",x"6C",x"66",x"66",x"66",x"66", -- 0x0440
    x"66",x"66",x"6C",x"F8",x"00",x"00",x"00",x"00", -- 0x0448
    x"00",x"00",x"FE",x"66",x"62",x"68",x"78",x"68", -- 0x0450
    x"60",x"62",x"66",x"FE",x"00",x"00",x"00",x"00", -- 0x0458
    x"00",x"00",x"FE",x"66",x"62",x"68",x"78",x"68", -- 0x0460
    x"60",x"60",x"60",x"F0",x"00",x"00",x"00",x"00", -- 0x0468
    x"00",x"00",x"3C",x"66",x"C2",x"C0",x"C0",x"DE", -- 0x0470
    x"C6",x"C6",x"66",x"3A",x"00",x"00",x"00",x"00", -- 0x0478
    x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"FE",x"C6", -- 0x0480
    x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x0488
    x"00",x"00",x"3C",x"18",x"18",x"18",x"18",x"18", -- 0x0490
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0498
    x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x04A0
    x"CC",x"CC",x"CC",x"78",x"00",x"00",x"00",x"00", -- 0x04A8
    x"00",x"00",x"E6",x"66",x"66",x"6C",x"78",x"78", -- 0x04B0
    x"6C",x"66",x"66",x"E6",x"00",x"00",x"00",x"00", -- 0x04B8
    x"00",x"00",x"F0",x"60",x"60",x"60",x"60",x"60", -- 0x04C0
    x"60",x"62",x"66",x"FE",x"00",x"00",x"00",x"00", -- 0x04C8
    x"00",x"00",x"C3",x"E7",x"FF",x"FF",x"DB",x"C3", -- 0x04D0
    x"C3",x"C3",x"C3",x"C3",x"00",x"00",x"00",x"00", -- 0x04D8
    x"00",x"00",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE", -- 0x04E0
    x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x04E8
    x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6", -- 0x04F0
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x04F8
    x"00",x"00",x"FC",x"66",x"66",x"66",x"7C",x"60", -- 0x0500
    x"60",x"60",x"60",x"F0",x"00",x"00",x"00",x"00", -- 0x0508
    x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6", -- 0x0510
    x"C6",x"D6",x"DE",x"7C",x"0C",x"0E",x"00",x"00", -- 0x0518
    x"00",x"00",x"FC",x"66",x"66",x"66",x"7C",x"6C", -- 0x0520
    x"66",x"66",x"66",x"E6",x"00",x"00",x"00",x"00", -- 0x0528
    x"00",x"00",x"7C",x"C6",x"C6",x"60",x"38",x"0C", -- 0x0530
    x"06",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0538
    x"00",x"00",x"FF",x"DB",x"99",x"18",x"18",x"18", -- 0x0540
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0548
    x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6", -- 0x0550
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0558
    x"00",x"00",x"C3",x"C3",x"C3",x"C3",x"C3",x"C3", -- 0x0560
    x"C3",x"66",x"3C",x"18",x"00",x"00",x"00",x"00", -- 0x0568
    x"00",x"00",x"C3",x"C3",x"C3",x"C3",x"C3",x"DB", -- 0x0570
    x"DB",x"FF",x"66",x"66",x"00",x"00",x"00",x"00", -- 0x0578
    x"00",x"00",x"C3",x"C3",x"66",x"3C",x"18",x"18", -- 0x0580
    x"3C",x"66",x"C3",x"C3",x"00",x"00",x"00",x"00", -- 0x0588
    x"00",x"00",x"C3",x"C3",x"C3",x"66",x"3C",x"18", -- 0x0590
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0598
    x"00",x"00",x"FF",x"C3",x"86",x"0C",x"18",x"30", -- 0x05A0
    x"60",x"C1",x"C3",x"FF",x"00",x"00",x"00",x"00", -- 0x05A8
    x"00",x"00",x"3C",x"30",x"30",x"30",x"30",x"30", -- 0x05B0
    x"30",x"30",x"30",x"3C",x"00",x"00",x"00",x"00", -- 0x05B8
    x"00",x"00",x"00",x"80",x"C0",x"E0",x"70",x"38", -- 0x05C0
    x"1C",x"0E",x"06",x"02",x"00",x"00",x"00",x"00", -- 0x05C8
    x"00",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x05D0
    x"0C",x"0C",x"0C",x"3C",x"00",x"00",x"00",x"00", -- 0x05D8
    x"10",x"38",x"6C",x"C6",x"00",x"00",x"00",x"00", -- 0x05E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F0
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00", -- 0x05F8
    x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00", -- 0x0600
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
    x"00",x"00",x"00",x"00",x"00",x"78",x"0C",x"7C", -- 0x0610
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0618
    x"00",x"00",x"E0",x"60",x"60",x"78",x"6C",x"66", -- 0x0620
    x"66",x"66",x"66",x"7C",x"00",x"00",x"00",x"00", -- 0x0628
    x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C0", -- 0x0630
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0638
    x"00",x"00",x"1C",x"0C",x"0C",x"3C",x"6C",x"CC", -- 0x0640
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0648
    x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"FE", -- 0x0650
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0658
    x"00",x"00",x"38",x"6C",x"64",x"60",x"F0",x"60", -- 0x0660
    x"60",x"60",x"60",x"F0",x"00",x"00",x"00",x"00", -- 0x0668
    x"00",x"00",x"00",x"00",x"00",x"76",x"CC",x"CC", -- 0x0670
    x"CC",x"CC",x"CC",x"7C",x"0C",x"CC",x"78",x"00", -- 0x0678
    x"00",x"00",x"E0",x"60",x"60",x"6C",x"76",x"66", -- 0x0680
    x"66",x"66",x"66",x"E6",x"00",x"00",x"00",x"00", -- 0x0688
    x"00",x"00",x"18",x"18",x"00",x"38",x"18",x"18", -- 0x0690
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0698
    x"00",x"00",x"06",x"06",x"00",x"0E",x"06",x"06", -- 0x06A0
    x"06",x"06",x"06",x"06",x"66",x"66",x"3C",x"00", -- 0x06A8
    x"00",x"00",x"E0",x"60",x"60",x"66",x"6C",x"78", -- 0x06B0
    x"78",x"6C",x"66",x"E6",x"00",x"00",x"00",x"00", -- 0x06B8
    x"00",x"00",x"38",x"18",x"18",x"18",x"18",x"18", -- 0x06C0
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x06C8
    x"00",x"00",x"00",x"00",x"00",x"E6",x"FF",x"DB", -- 0x06D0
    x"DB",x"DB",x"DB",x"DB",x"00",x"00",x"00",x"00", -- 0x06D8
    x"00",x"00",x"00",x"00",x"00",x"DC",x"66",x"66", -- 0x06E0
    x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"00", -- 0x06E8
    x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6", -- 0x06F0
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x06F8
    x"00",x"00",x"00",x"00",x"00",x"DC",x"66",x"66", -- 0x0700
    x"66",x"66",x"66",x"7C",x"60",x"60",x"F0",x"00", -- 0x0708
    x"00",x"00",x"00",x"00",x"00",x"76",x"CC",x"CC", -- 0x0710
    x"CC",x"CC",x"CC",x"7C",x"0C",x"0C",x"1E",x"00", -- 0x0718
    x"00",x"00",x"00",x"00",x"00",x"DC",x"76",x"66", -- 0x0720
    x"60",x"60",x"60",x"F0",x"00",x"00",x"00",x"00", -- 0x0728
    x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"60", -- 0x0730
    x"38",x"0C",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0738
    x"00",x"00",x"10",x"30",x"30",x"FC",x"30",x"30", -- 0x0740
    x"30",x"30",x"36",x"1C",x"00",x"00",x"00",x"00", -- 0x0748
    x"00",x"00",x"00",x"00",x"00",x"CC",x"CC",x"CC", -- 0x0750
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0758
    x"00",x"00",x"00",x"00",x"00",x"C3",x"C3",x"C3", -- 0x0760
    x"C3",x"66",x"3C",x"18",x"00",x"00",x"00",x"00", -- 0x0768
    x"00",x"00",x"00",x"00",x"00",x"C3",x"C3",x"C3", -- 0x0770
    x"DB",x"DB",x"FF",x"66",x"00",x"00",x"00",x"00", -- 0x0778
    x"00",x"00",x"00",x"00",x"00",x"C3",x"66",x"3C", -- 0x0780
    x"18",x"3C",x"66",x"C3",x"00",x"00",x"00",x"00", -- 0x0788
    x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6", -- 0x0790
    x"C6",x"C6",x"C6",x"7E",x"06",x"0C",x"F8",x"00", -- 0x0798
    x"00",x"00",x"00",x"00",x"00",x"FE",x"CC",x"18", -- 0x07A0
    x"30",x"60",x"C6",x"FE",x"00",x"00",x"00",x"00", -- 0x07A8
    x"00",x"00",x"0E",x"18",x"18",x"18",x"70",x"18", -- 0x07B0
    x"18",x"18",x"18",x"0E",x"00",x"00",x"00",x"00", -- 0x07B8
    x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"18", -- 0x07C0
    x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"00",x"70",x"18",x"18",x"18",x"0E",x"18", -- 0x07D0
    x"18",x"18",x"18",x"70",x"00",x"00",x"00",x"00", -- 0x07D8
    x"00",x"00",x"76",x"DC",x"00",x"00",x"00",x"00", -- 0x07E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
    x"00",x"00",x"00",x"00",x"10",x"38",x"6C",x"C6", -- 0x07F0
    x"C6",x"C6",x"FE",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
    x"00",x"00",x"3C",x"66",x"C2",x"C0",x"C0",x"C0", -- 0x0800
    x"C2",x"66",x"3C",x"0C",x"06",x"7C",x"00",x"00", -- 0x0808
    x"00",x"00",x"CC",x"00",x"00",x"CC",x"CC",x"CC", -- 0x0810
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0818
    x"00",x"0C",x"18",x"30",x"00",x"7C",x"C6",x"FE", -- 0x0820
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0828
    x"00",x"10",x"38",x"6C",x"00",x"78",x"0C",x"7C", -- 0x0830
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0838
    x"00",x"00",x"CC",x"00",x"00",x"78",x"0C",x"7C", -- 0x0840
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0848
    x"00",x"60",x"30",x"18",x"00",x"78",x"0C",x"7C", -- 0x0850
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0858
    x"00",x"38",x"6C",x"38",x"00",x"78",x"0C",x"7C", -- 0x0860
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0868
    x"00",x"00",x"00",x"00",x"3C",x"66",x"60",x"60", -- 0x0870
    x"66",x"3C",x"0C",x"06",x"3C",x"00",x"00",x"00", -- 0x0878
    x"00",x"10",x"38",x"6C",x"00",x"7C",x"C6",x"FE", -- 0x0880
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0888
    x"00",x"00",x"C6",x"00",x"00",x"7C",x"C6",x"FE", -- 0x0890
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0898
    x"00",x"60",x"30",x"18",x"00",x"7C",x"C6",x"FE", -- 0x08A0
    x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x08A8
    x"00",x"00",x"66",x"00",x"00",x"38",x"18",x"18", -- 0x08B0
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x08B8
    x"00",x"18",x"3C",x"66",x"00",x"38",x"18",x"18", -- 0x08C0
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x08C8
    x"00",x"60",x"30",x"18",x"00",x"38",x"18",x"18", -- 0x08D0
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x08D8
    x"00",x"C6",x"00",x"10",x"38",x"6C",x"C6",x"C6", -- 0x08E0
    x"FE",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x08E8
    x"38",x"6C",x"38",x"00",x"38",x"6C",x"C6",x"C6", -- 0x08F0
    x"FE",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x08F8
    x"18",x"30",x"60",x"00",x"FE",x"66",x"60",x"7C", -- 0x0900
    x"60",x"60",x"66",x"FE",x"00",x"00",x"00",x"00", -- 0x0908
    x"00",x"00",x"00",x"00",x"00",x"6E",x"3B",x"1B", -- 0x0910
    x"7E",x"D8",x"DC",x"77",x"00",x"00",x"00",x"00", -- 0x0918
    x"00",x"00",x"3E",x"6C",x"CC",x"CC",x"FE",x"CC", -- 0x0920
    x"CC",x"CC",x"CC",x"CE",x"00",x"00",x"00",x"00", -- 0x0928
    x"00",x"10",x"38",x"6C",x"00",x"7C",x"C6",x"C6", -- 0x0930
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0938
    x"00",x"00",x"C6",x"00",x"00",x"7C",x"C6",x"C6", -- 0x0940
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0948
    x"00",x"60",x"30",x"18",x"00",x"7C",x"C6",x"C6", -- 0x0950
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0958
    x"00",x"30",x"78",x"CC",x"00",x"CC",x"CC",x"CC", -- 0x0960
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0968
    x"00",x"60",x"30",x"18",x"00",x"CC",x"CC",x"CC", -- 0x0970
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0978
    x"00",x"00",x"C6",x"00",x"00",x"C6",x"C6",x"C6", -- 0x0980
    x"C6",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00", -- 0x0988
    x"00",x"C6",x"00",x"7C",x"C6",x"C6",x"C6",x"C6", -- 0x0990
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0998
    x"00",x"C6",x"00",x"C6",x"C6",x"C6",x"C6",x"C6", -- 0x09A0
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x09A8
    x"00",x"18",x"18",x"7E",x"C3",x"C0",x"C0",x"C0", -- 0x09B0
    x"C3",x"7E",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x09B8
    x"00",x"38",x"6C",x"64",x"60",x"F0",x"60",x"60", -- 0x09C0
    x"60",x"60",x"E6",x"FC",x"00",x"00",x"00",x"00", -- 0x09C8
    x"00",x"00",x"C3",x"66",x"3C",x"18",x"FF",x"18", -- 0x09D0
    x"FF",x"18",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x09D8
    x"00",x"FC",x"66",x"66",x"7C",x"62",x"66",x"6F", -- 0x09E0
    x"66",x"66",x"66",x"F3",x"00",x"00",x"00",x"00", -- 0x09E8
    x"00",x"0E",x"1B",x"18",x"18",x"18",x"7E",x"18", -- 0x09F0
    x"18",x"18",x"18",x"18",x"D8",x"70",x"00",x"00", -- 0x09F8
    x"00",x"18",x"30",x"60",x"00",x"78",x"0C",x"7C", -- 0x0A00
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0A08
    x"00",x"0C",x"18",x"30",x"00",x"38",x"18",x"18", -- 0x0A10
    x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00", -- 0x0A18
    x"00",x"18",x"30",x"60",x"00",x"7C",x"C6",x"C6", -- 0x0A20
    x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0A28
    x"00",x"18",x"30",x"60",x"00",x"CC",x"CC",x"CC", -- 0x0A30
    x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",x"00", -- 0x0A38
    x"00",x"00",x"76",x"DC",x"00",x"DC",x"66",x"66", -- 0x0A40
    x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"00", -- 0x0A48
    x"76",x"DC",x"00",x"C6",x"E6",x"F6",x"FE",x"DE", -- 0x0A50
    x"CE",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x0A58
    x"00",x"3C",x"6C",x"6C",x"3E",x"00",x"7E",x"00", -- 0x0A60
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A68
    x"00",x"38",x"6C",x"6C",x"38",x"00",x"7C",x"00", -- 0x0A70
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A78
    x"00",x"00",x"30",x"30",x"00",x"30",x"30",x"60", -- 0x0A80
    x"C0",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00", -- 0x0A88
    x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"C0", -- 0x0A90
    x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x0A98
    x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"06", -- 0x0AA0
    x"06",x"06",x"06",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
    x"00",x"C0",x"C0",x"C2",x"C6",x"CC",x"18",x"30", -- 0x0AB0
    x"60",x"CE",x"9B",x"06",x"0C",x"1F",x"00",x"00", -- 0x0AB8
    x"00",x"C0",x"C0",x"C2",x"C6",x"CC",x"18",x"30", -- 0x0AC0
    x"66",x"CE",x"96",x"3E",x"06",x"06",x"00",x"00", -- 0x0AC8
    x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"18", -- 0x0AD0
    x"3C",x"3C",x"3C",x"18",x"00",x"00",x"00",x"00", -- 0x0AD8
    x"00",x"00",x"00",x"00",x"00",x"36",x"6C",x"D8", -- 0x0AE0
    x"6C",x"36",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE8
    x"00",x"00",x"00",x"00",x"00",x"D8",x"6C",x"36", -- 0x0AF0
    x"6C",x"D8",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF8
    x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44", -- 0x0B00
    x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44", -- 0x0B08
    x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA", -- 0x0B10
    x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA", -- 0x0B18
    x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77", -- 0x0B20
    x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77", -- 0x0B28
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0B30
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0B38
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"F8", -- 0x0B40
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0B48
    x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"F8", -- 0x0B50
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0B58
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"F6", -- 0x0B60
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0B68
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE", -- 0x0B70
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0B78
    x"00",x"00",x"00",x"00",x"00",x"F8",x"18",x"F8", -- 0x0B80
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0B88
    x"36",x"36",x"36",x"36",x"36",x"F6",x"06",x"F6", -- 0x0B90
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0B98
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0BA0
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0BA8
    x"00",x"00",x"00",x"00",x"00",x"FE",x"06",x"F6", -- 0x0BB0
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0BB8
    x"36",x"36",x"36",x"36",x"36",x"F6",x"06",x"FE", -- 0x0BC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC8
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FE", -- 0x0BD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD8
    x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"F8", -- 0x0BE0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8", -- 0x0BF0
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0BF8
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F", -- 0x0C00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C08
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"FF", -- 0x0C10
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x0C20
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0C28
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F", -- 0x0C30
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0C38
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x0C40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C48
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"FF", -- 0x0C50
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0C58
    x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"1F", -- 0x0C60
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0C68
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37", -- 0x0C70
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0C78
    x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"3F", -- 0x0C80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C88
    x"00",x"00",x"00",x"00",x"00",x"3F",x"30",x"37", -- 0x0C90
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0C98
    x"36",x"36",x"36",x"36",x"36",x"F7",x"00",x"FF", -- 0x0CA0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"F7", -- 0x0CB0
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0CB8
    x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"37", -- 0x0CC0
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0CC8
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF", -- 0x0CD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD8
    x"36",x"36",x"36",x"36",x"36",x"F7",x"00",x"F7", -- 0x0CE0
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0CE8
    x"18",x"18",x"18",x"18",x"18",x"FF",x"00",x"FF", -- 0x0CF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FF", -- 0x0D00
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D08
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF", -- 0x0D10
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0D18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x0D20
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0D28
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3F", -- 0x0D30
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D38
    x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"1F", -- 0x0D40
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D48
    x"00",x"00",x"00",x"00",x"00",x"1F",x"18",x"1F", -- 0x0D50
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0D58
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F", -- 0x0D60
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0D68
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FF", -- 0x0D70
    x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36", -- 0x0D78
    x"18",x"18",x"18",x"18",x"18",x"FF",x"18",x"FF", -- 0x0D80
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0D88
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"F8", -- 0x0D90
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F", -- 0x0DA0
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x0DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC8
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0DD0
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0DD8
    x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0DE0
    x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0DE8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x0DF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF8
    x"00",x"00",x"00",x"00",x"00",x"76",x"DC",x"D8", -- 0x0E00
    x"D8",x"D8",x"DC",x"76",x"00",x"00",x"00",x"00", -- 0x0E08
    x"00",x"00",x"78",x"CC",x"CC",x"CC",x"D8",x"CC", -- 0x0E10
    x"C6",x"C6",x"C6",x"CC",x"00",x"00",x"00",x"00", -- 0x0E18
    x"00",x"00",x"FE",x"C6",x"C6",x"C0",x"C0",x"C0", -- 0x0E20
    x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00", -- 0x0E28
    x"00",x"00",x"00",x"00",x"FE",x"6C",x"6C",x"6C", -- 0x0E30
    x"6C",x"6C",x"6C",x"6C",x"00",x"00",x"00",x"00", -- 0x0E38
    x"00",x"00",x"00",x"FE",x"C6",x"60",x"30",x"18", -- 0x0E40
    x"30",x"60",x"C6",x"FE",x"00",x"00",x"00",x"00", -- 0x0E48
    x"00",x"00",x"00",x"00",x"00",x"7E",x"D8",x"D8", -- 0x0E50
    x"D8",x"D8",x"D8",x"70",x"00",x"00",x"00",x"00", -- 0x0E58
    x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"66", -- 0x0E60
    x"66",x"7C",x"60",x"60",x"C0",x"00",x"00",x"00", -- 0x0E68
    x"00",x"00",x"00",x"00",x"76",x"DC",x"18",x"18", -- 0x0E70
    x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00", -- 0x0E78
    x"00",x"00",x"00",x"7E",x"18",x"3C",x"66",x"66", -- 0x0E80
    x"66",x"3C",x"18",x"7E",x"00",x"00",x"00",x"00", -- 0x0E88
    x"00",x"00",x"00",x"38",x"6C",x"C6",x"C6",x"FE", -- 0x0E90
    x"C6",x"C6",x"6C",x"38",x"00",x"00",x"00",x"00", -- 0x0E98
    x"00",x"00",x"38",x"6C",x"C6",x"C6",x"C6",x"6C", -- 0x0EA0
    x"6C",x"6C",x"6C",x"EE",x"00",x"00",x"00",x"00", -- 0x0EA8
    x"00",x"00",x"1E",x"30",x"18",x"0C",x"3E",x"66", -- 0x0EB0
    x"66",x"66",x"66",x"3C",x"00",x"00",x"00",x"00", -- 0x0EB8
    x"00",x"00",x"00",x"00",x"00",x"7E",x"DB",x"DB", -- 0x0EC0
    x"DB",x"7E",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC8
    x"00",x"00",x"00",x"03",x"06",x"7E",x"DB",x"DB", -- 0x0ED0
    x"F3",x"7E",x"60",x"C0",x"00",x"00",x"00",x"00", -- 0x0ED8
    x"00",x"00",x"1C",x"30",x"60",x"60",x"7C",x"60", -- 0x0EE0
    x"60",x"60",x"30",x"1C",x"00",x"00",x"00",x"00", -- 0x0EE8
    x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6", -- 0x0EF0
    x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"FE", -- 0x0F00
    x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00", -- 0x0F08
    x"00",x"00",x"00",x"00",x"18",x"18",x"7E",x"18", -- 0x0F10
    x"18",x"00",x"00",x"FF",x"00",x"00",x"00",x"00", -- 0x0F18
    x"00",x"00",x"00",x"30",x"18",x"0C",x"06",x"0C", -- 0x0F20
    x"18",x"30",x"00",x"7E",x"00",x"00",x"00",x"00", -- 0x0F28
    x"00",x"00",x"00",x"0C",x"18",x"30",x"60",x"30", -- 0x0F30
    x"18",x"0C",x"00",x"7E",x"00",x"00",x"00",x"00", -- 0x0F38
    x"00",x"00",x"0E",x"1B",x"1B",x"1B",x"18",x"18", -- 0x0F40
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0F48
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- 0x0F50
    x"D8",x"D8",x"D8",x"70",x"00",x"00",x"00",x"00", -- 0x0F58
    x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"7E", -- 0x0F60
    x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00", -- 0x0F68
    x"00",x"00",x"00",x"00",x"00",x"76",x"DC",x"00", -- 0x0F70
    x"76",x"DC",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F78
    x"00",x"38",x"6C",x"6C",x"38",x"00",x"00",x"00", -- 0x0F80
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F88
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- 0x0F90
    x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F98
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA0
    x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA8
    x"00",x"0F",x"0C",x"0C",x"0C",x"0C",x"0C",x"EC", -- 0x0FB0
    x"6C",x"6C",x"3C",x"1C",x"00",x"00",x"00",x"00", -- 0x0FB8
    x"00",x"D8",x"6C",x"6C",x"6C",x"6C",x"6C",x"00", -- 0x0FC0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC8
    x"00",x"70",x"D8",x"30",x"60",x"C8",x"F8",x"00", -- 0x0FD0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
    x"00",x"00",x"00",x"00",x"7C",x"7C",x"7C",x"7C", -- 0x0FE0
    x"7C",x"7C",x"7C",x"00",x"00",x"00",x"00",x"00", -- 0x0FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
